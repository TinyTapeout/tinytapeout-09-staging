module tt_um_kmakise_sram (clk,
    ena,
    rst_n,
    VDPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VDPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \SRAMController_ins.addr[0] ;
 wire \SRAMController_ins.addr[1] ;
 wire \SRAMController_ins.addr[2] ;
 wire \SRAMController_ins.addr[3] ;
 wire \SRAMController_ins.addr_tmp[0] ;
 wire \SRAMController_ins.addr_tmp[1] ;
 wire \SRAMController_ins.addr_tmp[2] ;
 wire \SRAMController_ins.addr_tmp[3] ;
 wire \SRAMController_ins.csb_n ;
 wire \SRAMController_ins.cur_state[0] ;
 wire \SRAMController_ins.cur_state[1] ;
 wire \SRAMController_ins.cur_state[2] ;
 wire \SRAMController_ins.cur_state[3] ;
 wire \SRAMController_ins.data_tmp[0] ;
 wire \SRAMController_ins.data_tmp[10] ;
 wire \SRAMController_ins.data_tmp[11] ;
 wire \SRAMController_ins.data_tmp[12] ;
 wire \SRAMController_ins.data_tmp[13] ;
 wire \SRAMController_ins.data_tmp[14] ;
 wire \SRAMController_ins.data_tmp[15] ;
 wire \SRAMController_ins.data_tmp[16] ;
 wire \SRAMController_ins.data_tmp[17] ;
 wire \SRAMController_ins.data_tmp[18] ;
 wire \SRAMController_ins.data_tmp[19] ;
 wire \SRAMController_ins.data_tmp[1] ;
 wire \SRAMController_ins.data_tmp[20] ;
 wire \SRAMController_ins.data_tmp[21] ;
 wire \SRAMController_ins.data_tmp[22] ;
 wire \SRAMController_ins.data_tmp[23] ;
 wire \SRAMController_ins.data_tmp[24] ;
 wire \SRAMController_ins.data_tmp[25] ;
 wire \SRAMController_ins.data_tmp[26] ;
 wire \SRAMController_ins.data_tmp[27] ;
 wire \SRAMController_ins.data_tmp[28] ;
 wire \SRAMController_ins.data_tmp[29] ;
 wire \SRAMController_ins.data_tmp[2] ;
 wire \SRAMController_ins.data_tmp[30] ;
 wire \SRAMController_ins.data_tmp[31] ;
 wire \SRAMController_ins.data_tmp[3] ;
 wire \SRAMController_ins.data_tmp[4] ;
 wire \SRAMController_ins.data_tmp[5] ;
 wire \SRAMController_ins.data_tmp[6] ;
 wire \SRAMController_ins.data_tmp[7] ;
 wire \SRAMController_ins.data_tmp[8] ;
 wire \SRAMController_ins.data_tmp[9] ;
 wire \SRAMController_ins.nxt_state[0] ;
 wire \SRAMController_ins.nxt_state[1] ;
 wire \SRAMController_ins.nxt_state[2] ;
 wire \SRAMController_ins.nxt_state[3] ;
 wire \SRAMController_ins.rx_data_out[0] ;
 wire \SRAMController_ins.rx_data_out[1] ;
 wire \SRAMController_ins.rx_data_out[2] ;
 wire \SRAMController_ins.rx_data_out[3] ;
 wire \SRAMController_ins.rx_data_out[4] ;
 wire \SRAMController_ins.rx_data_out[5] ;
 wire \SRAMController_ins.rx_data_out[6] ;
 wire \SRAMController_ins.rx_data_out[7] ;
 wire \SRAMController_ins.rx_valid ;
 wire \SRAMController_ins.sram_data_in[0] ;
 wire \SRAMController_ins.sram_data_in[10] ;
 wire \SRAMController_ins.sram_data_in[11] ;
 wire \SRAMController_ins.sram_data_in[12] ;
 wire \SRAMController_ins.sram_data_in[13] ;
 wire \SRAMController_ins.sram_data_in[14] ;
 wire \SRAMController_ins.sram_data_in[15] ;
 wire \SRAMController_ins.sram_data_in[16] ;
 wire \SRAMController_ins.sram_data_in[17] ;
 wire \SRAMController_ins.sram_data_in[18] ;
 wire \SRAMController_ins.sram_data_in[19] ;
 wire \SRAMController_ins.sram_data_in[1] ;
 wire \SRAMController_ins.sram_data_in[20] ;
 wire \SRAMController_ins.sram_data_in[21] ;
 wire \SRAMController_ins.sram_data_in[22] ;
 wire \SRAMController_ins.sram_data_in[23] ;
 wire \SRAMController_ins.sram_data_in[24] ;
 wire \SRAMController_ins.sram_data_in[25] ;
 wire \SRAMController_ins.sram_data_in[26] ;
 wire \SRAMController_ins.sram_data_in[27] ;
 wire \SRAMController_ins.sram_data_in[28] ;
 wire \SRAMController_ins.sram_data_in[29] ;
 wire \SRAMController_ins.sram_data_in[2] ;
 wire \SRAMController_ins.sram_data_in[30] ;
 wire \SRAMController_ins.sram_data_in[31] ;
 wire \SRAMController_ins.sram_data_in[3] ;
 wire \SRAMController_ins.sram_data_in[4] ;
 wire \SRAMController_ins.sram_data_in[5] ;
 wire \SRAMController_ins.sram_data_in[6] ;
 wire \SRAMController_ins.sram_data_in[7] ;
 wire \SRAMController_ins.sram_data_in[8] ;
 wire \SRAMController_ins.sram_data_in[9] ;
 wire \SRAMController_ins.sram_data_out[0] ;
 wire \SRAMController_ins.sram_data_out[10] ;
 wire \SRAMController_ins.sram_data_out[11] ;
 wire \SRAMController_ins.sram_data_out[12] ;
 wire \SRAMController_ins.sram_data_out[13] ;
 wire \SRAMController_ins.sram_data_out[14] ;
 wire \SRAMController_ins.sram_data_out[15] ;
 wire \SRAMController_ins.sram_data_out[16] ;
 wire \SRAMController_ins.sram_data_out[17] ;
 wire \SRAMController_ins.sram_data_out[18] ;
 wire \SRAMController_ins.sram_data_out[19] ;
 wire \SRAMController_ins.sram_data_out[1] ;
 wire \SRAMController_ins.sram_data_out[20] ;
 wire \SRAMController_ins.sram_data_out[21] ;
 wire \SRAMController_ins.sram_data_out[22] ;
 wire \SRAMController_ins.sram_data_out[23] ;
 wire \SRAMController_ins.sram_data_out[24] ;
 wire \SRAMController_ins.sram_data_out[25] ;
 wire \SRAMController_ins.sram_data_out[26] ;
 wire \SRAMController_ins.sram_data_out[27] ;
 wire \SRAMController_ins.sram_data_out[28] ;
 wire \SRAMController_ins.sram_data_out[29] ;
 wire \SRAMController_ins.sram_data_out[2] ;
 wire \SRAMController_ins.sram_data_out[30] ;
 wire \SRAMController_ins.sram_data_out[31] ;
 wire \SRAMController_ins.sram_data_out[3] ;
 wire \SRAMController_ins.sram_data_out[4] ;
 wire \SRAMController_ins.sram_data_out[5] ;
 wire \SRAMController_ins.sram_data_out[6] ;
 wire \SRAMController_ins.sram_data_out[7] ;
 wire \SRAMController_ins.sram_data_out[8] ;
 wire \SRAMController_ins.sram_data_out[9] ;
 wire \SRAMController_ins.sram_tmp[0] ;
 wire \SRAMController_ins.sram_tmp[10] ;
 wire \SRAMController_ins.sram_tmp[11] ;
 wire \SRAMController_ins.sram_tmp[12] ;
 wire \SRAMController_ins.sram_tmp[13] ;
 wire \SRAMController_ins.sram_tmp[14] ;
 wire \SRAMController_ins.sram_tmp[15] ;
 wire \SRAMController_ins.sram_tmp[16] ;
 wire \SRAMController_ins.sram_tmp[17] ;
 wire \SRAMController_ins.sram_tmp[18] ;
 wire \SRAMController_ins.sram_tmp[19] ;
 wire \SRAMController_ins.sram_tmp[1] ;
 wire \SRAMController_ins.sram_tmp[20] ;
 wire \SRAMController_ins.sram_tmp[21] ;
 wire \SRAMController_ins.sram_tmp[22] ;
 wire \SRAMController_ins.sram_tmp[23] ;
 wire \SRAMController_ins.sram_tmp[24] ;
 wire \SRAMController_ins.sram_tmp[25] ;
 wire \SRAMController_ins.sram_tmp[26] ;
 wire \SRAMController_ins.sram_tmp[27] ;
 wire \SRAMController_ins.sram_tmp[28] ;
 wire \SRAMController_ins.sram_tmp[29] ;
 wire \SRAMController_ins.sram_tmp[2] ;
 wire \SRAMController_ins.sram_tmp[30] ;
 wire \SRAMController_ins.sram_tmp[31] ;
 wire \SRAMController_ins.sram_tmp[3] ;
 wire \SRAMController_ins.sram_tmp[4] ;
 wire \SRAMController_ins.sram_tmp[5] ;
 wire \SRAMController_ins.sram_tmp[6] ;
 wire \SRAMController_ins.sram_tmp[7] ;
 wire \SRAMController_ins.sram_tmp[8] ;
 wire \SRAMController_ins.sram_tmp[9] ;
 wire \SRAMController_ins.tx_ready ;
 wire \SRAMController_ins.we_n ;
 wire \UARTReceiver_ins.bitIndex[0] ;
 wire \UARTReceiver_ins.bitIndex[1] ;
 wire \UARTReceiver_ins.bitIndex[2] ;
 wire \UARTReceiver_ins.data[0] ;
 wire \UARTReceiver_ins.data[1] ;
 wire \UARTReceiver_ins.data[2] ;
 wire \UARTReceiver_ins.data[3] ;
 wire \UARTReceiver_ins.data[4] ;
 wire \UARTReceiver_ins.data[5] ;
 wire \UARTReceiver_ins.data[6] ;
 wire \UARTReceiver_ins.data[7] ;
 wire \UARTReceiver_ins.error ;
 wire \UARTReceiver_ins.inputReg[0] ;
 wire \UARTReceiver_ins.inputReg[1] ;
 wire \UARTReceiver_ins.inputReg[2] ;
 wire \UARTReceiver_ins.out_latched ;
 wire \UARTReceiver_ins.overrun ;
 wire \UARTReceiver_ins.rxCounter[0] ;
 wire \UARTReceiver_ins.rxCounter[1] ;
 wire \UARTReceiver_ins.rxCounter[2] ;
 wire \UARTReceiver_ins.rxCounter[3] ;
 wire \UARTReceiver_ins.rxCounter[4] ;
 wire \UARTReceiver_ins.rxCounter[5] ;
 wire \UARTReceiver_ins.rxCounter[6] ;
 wire \UARTReceiver_ins.rxCounter[7] ;
 wire \UARTReceiver_ins.sampleCount[0] ;
 wire \UARTReceiver_ins.sampleCount[1] ;
 wire \UARTReceiver_ins.sampleCount[2] ;
 wire \UARTReceiver_ins.sampleCount[3] ;
 wire \UARTReceiver_ins.state[0] ;
 wire \UARTReceiver_ins.state[1] ;
 wire \UARTReceiver_ins.state[2] ;
 wire \UARTReceiver_ins.state[3] ;
 wire \UARTTransmitter_ins.bitIndex[0] ;
 wire \UARTTransmitter_ins.bitIndex[1] ;
 wire \UARTTransmitter_ins.bitIndex[2] ;
 wire \UARTTransmitter_ins.data[0] ;
 wire \UARTTransmitter_ins.data[1] ;
 wire \UARTTransmitter_ins.data[2] ;
 wire \UARTTransmitter_ins.data[3] ;
 wire \UARTTransmitter_ins.data[4] ;
 wire \UARTTransmitter_ins.data[5] ;
 wire \UARTTransmitter_ins.data[6] ;
 wire \UARTTransmitter_ins.data[7] ;
 wire \UARTTransmitter_ins.out ;
 wire \UARTTransmitter_ins.state[0] ;
 wire \UARTTransmitter_ins.state[1] ;
 wire \UARTTransmitter_ins.state[2] ;
 wire \UARTTransmitter_ins.state[3] ;
 wire \UARTTransmitter_ins.txCounter[0] ;
 wire \UARTTransmitter_ins.txCounter[10] ;
 wire \UARTTransmitter_ins.txCounter[11] ;
 wire \UARTTransmitter_ins.txCounter[1] ;
 wire \UARTTransmitter_ins.txCounter[2] ;
 wire \UARTTransmitter_ins.txCounter[3] ;
 wire \UARTTransmitter_ins.txCounter[4] ;
 wire \UARTTransmitter_ins.txCounter[5] ;
 wire \UARTTransmitter_ins.txCounter[6] ;
 wire \UARTTransmitter_ins.txCounter[7] ;
 wire \UARTTransmitter_ins.txCounter[8] ;
 wire \UARTTransmitter_ins.txCounter[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire net56;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire clknet_0_clk;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;

 sky130_fd_sc_hd__or2_1 _0518_ (.A(\UARTReceiver_ins.rxCounter[0] ),
    .B(\UARTReceiver_ins.rxCounter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0139_));
 sky130_fd_sc_hd__o41a_4 _0519_ (.A1(\UARTReceiver_ins.rxCounter[4] ),
    .A2(\UARTReceiver_ins.rxCounter[3] ),
    .A3(\UARTReceiver_ins.rxCounter[2] ),
    .A4(_0139_),
    .B1(\UARTReceiver_ins.rxCounter[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0140_));
 sky130_fd_sc_hd__o211ai_4 _0520_ (.A1(\UARTReceiver_ins.rxCounter[6] ),
    .A2(_0140_),
    .B1(net21),
    .C1(\UARTReceiver_ins.rxCounter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0141_));
 sky130_fd_sc_hd__nand3_1 _0521_ (.A(\UARTReceiver_ins.inputReg[2] ),
    .B(\UARTReceiver_ins.inputReg[1] ),
    .C(\UARTReceiver_ins.inputReg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0142_));
 sky130_fd_sc_hd__and4_1 _0522_ (.A(\UARTReceiver_ins.sampleCount[3] ),
    .B(\UARTReceiver_ins.sampleCount[2] ),
    .C(\UARTReceiver_ins.sampleCount[1] ),
    .D(\UARTReceiver_ins.sampleCount[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0143_));
 sky130_fd_sc_hd__and3_1 _0523_ (.A(net8),
    .B(_0142_),
    .C(_0143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0144_));
 sky130_fd_sc_hd__or3_1 _0524_ (.A(\UARTReceiver_ins.sampleCount[3] ),
    .B(\UARTReceiver_ins.sampleCount[1] ),
    .C(\UARTReceiver_ins.sampleCount[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0145_));
 sky130_fd_sc_hd__or2_1 _0525_ (.A(\UARTReceiver_ins.sampleCount[3] ),
    .B(\UARTReceiver_ins.sampleCount[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0146_));
 sky130_fd_sc_hd__inv_2 _0526_ (.A(\UARTReceiver_ins.state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0147_));
 sky130_fd_sc_hd__a21o_2 _0527_ (.A1(_0145_),
    .A2(_0146_),
    .B1(_0147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0148_));
 sky130_fd_sc_hd__or3_1 _0528_ (.A(\UARTReceiver_ins.inputReg[2] ),
    .B(\UARTReceiver_ins.inputReg[1] ),
    .C(\UARTReceiver_ins.inputReg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0149_));
 sky130_fd_sc_hd__o21ai_1 _0529_ (.A1(\UARTReceiver_ins.sampleCount[2] ),
    .A2(_0145_),
    .B1(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0150_));
 sky130_fd_sc_hd__nor2_1 _0530_ (.A(_0148_),
    .B(_0150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0151_));
 sky130_fd_sc_hd__o21ai_4 _0531_ (.A1(\UARTReceiver_ins.rxCounter[6] ),
    .A2(_0140_),
    .B1(\UARTReceiver_ins.rxCounter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0152_));
 sky130_fd_sc_hd__nand2_2 _0532_ (.A(net21),
    .B(_0152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0153_));
 sky130_fd_sc_hd__o32a_1 _0533_ (.A1(_0141_),
    .A2(_0144_),
    .A3(_0151_),
    .B1(_0153_),
    .B2(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0000_));
 sky130_fd_sc_hd__o21a_1 _0534_ (.A1(\UARTReceiver_ins.rxCounter[6] ),
    .A2(_0140_),
    .B1(\UARTReceiver_ins.rxCounter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0154_));
 sky130_fd_sc_hd__buf_2 _0535_ (.A(_0154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0155_));
 sky130_fd_sc_hd__and3_1 _0536_ (.A(\UARTReceiver_ins.bitIndex[2] ),
    .B(\UARTReceiver_ins.bitIndex[1] ),
    .C(\UARTReceiver_ins.bitIndex[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0156_));
 sky130_fd_sc_hd__and3_1 _0537_ (.A(_0155_),
    .B(_0143_),
    .C(_0156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0157_));
 sky130_fd_sc_hd__nand2_1 _0538_ (.A(net19),
    .B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0158_));
 sky130_fd_sc_hd__and3_1 _0539_ (.A(\UARTReceiver_ins.state[2] ),
    .B(_0145_),
    .C(_0146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _0540_ (.A(net19),
    .B(_0155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0160_));
 sky130_fd_sc_hd__a2bb2o_1 _0541_ (.A1_N(_0157_),
    .A2_N(_0158_),
    .B1(_0159_),
    .B2(_0160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0001_));
 sky130_fd_sc_hd__a21o_1 _0542_ (.A1(\UARTTransmitter_ins.txCounter[1] ),
    .A2(\UARTTransmitter_ins.txCounter[0] ),
    .B1(\UARTTransmitter_ins.txCounter[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0161_));
 sky130_fd_sc_hd__or4_1 _0543_ (.A(\UARTTransmitter_ins.txCounter[10] ),
    .B(\UARTTransmitter_ins.txCounter[8] ),
    .C(\UARTTransmitter_ins.txCounter[7] ),
    .D(\UARTTransmitter_ins.txCounter[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0162_));
 sky130_fd_sc_hd__and2_1 _0544_ (.A(\UARTTransmitter_ins.txCounter[5] ),
    .B(\UARTTransmitter_ins.txCounter[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0163_));
 sky130_fd_sc_hd__a311o_4 _0545_ (.A1(\UARTTransmitter_ins.txCounter[5] ),
    .A2(\UARTTransmitter_ins.txCounter[3] ),
    .A3(_0161_),
    .B1(_0162_),
    .C1(_0163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0164_));
 sky130_fd_sc_hd__o21a_2 _0546_ (.A1(\UARTTransmitter_ins.txCounter[10] ),
    .A2(\UARTTransmitter_ins.txCounter[9] ),
    .B1(\UARTTransmitter_ins.txCounter[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0165_));
 sky130_fd_sc_hd__nor4b_1 _0547_ (.A(\SRAMController_ins.cur_state[0] ),
    .B(\SRAMController_ins.cur_state[2] ),
    .C(\SRAMController_ins.cur_state[3] ),
    .D_N(\SRAMController_ins.cur_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0166_));
 sky130_fd_sc_hd__nor4b_1 _0548_ (.A(\SRAMController_ins.cur_state[1] ),
    .B(\SRAMController_ins.cur_state[0] ),
    .C(\SRAMController_ins.cur_state[3] ),
    .D_N(\SRAMController_ins.cur_state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0167_));
 sky130_fd_sc_hd__and4bb_1 _0549_ (.A_N(\SRAMController_ins.cur_state[1] ),
    .B_N(\SRAMController_ins.cur_state[3] ),
    .C(\SRAMController_ins.cur_state[2] ),
    .D(\SRAMController_ins.cur_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0168_));
 sky130_fd_sc_hd__and4bb_1 _0550_ (.A_N(\SRAMController_ins.cur_state[2] ),
    .B_N(\SRAMController_ins.cur_state[3] ),
    .C(\SRAMController_ins.cur_state[1] ),
    .D(\SRAMController_ins.cur_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0169_));
 sky130_fd_sc_hd__o41a_1 _0551_ (.A1(_0166_),
    .A2(_0167_),
    .A3(_0168_),
    .A4(_0169_),
    .B1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_4 _0552_ (.A(_0170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0171_));
 sky130_fd_sc_hd__a21oi_4 _0553_ (.A1(_0164_),
    .A2(_0165_),
    .B1(_0171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0172_));
 sky130_fd_sc_hd__clkbuf_8 _0554_ (.A(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0173_));
 sky130_fd_sc_hd__clkbuf_8 _0555_ (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0174_));
 sky130_fd_sc_hd__clkbuf_8 _0556_ (.A(_0168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0175_));
 sky130_fd_sc_hd__o41ai_1 _0557_ (.A1(_0173_),
    .A2(_0174_),
    .A3(_0175_),
    .A4(_0169_),
    .B1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0176_));
 sky130_fd_sc_hd__and4_1 _0558_ (.A(\UARTTransmitter_ins.state[1] ),
    .B(_0164_),
    .C(_0165_),
    .D(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0177_));
 sky130_fd_sc_hd__and3_1 _0559_ (.A(\UARTTransmitter_ins.bitIndex[2] ),
    .B(\UARTTransmitter_ins.bitIndex[1] ),
    .C(\UARTTransmitter_ins.bitIndex[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0178_));
 sky130_fd_sc_hd__a22o_1 _0560_ (.A1(\UARTTransmitter_ins.state[3] ),
    .A2(_0172_),
    .B1(_0177_),
    .B2(_0178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0179_));
 sky130_fd_sc_hd__and2_1 _0561_ (.A(net24),
    .B(_0179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0180_));
 sky130_fd_sc_hd__clkbuf_1 _0562_ (.A(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0007_));
 sky130_fd_sc_hd__and3_1 _0563_ (.A(_0164_),
    .B(_0165_),
    .C(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0181_));
 sky130_fd_sc_hd__nor2b_2 _0564_ (.A(_0181_),
    .B_N(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0182_));
 sky130_fd_sc_hd__o21a_1 _0565_ (.A1(net59),
    .A2(_0171_),
    .B1(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0006_));
 sky130_fd_sc_hd__nand2_1 _0566_ (.A(_0164_),
    .B(_0165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _0567_ (.A(_0178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0184_));
 sky130_fd_sc_hd__o2111a_1 _0568_ (.A1(_0183_),
    .A2(_0184_),
    .B1(net3),
    .C1(net24),
    .D1(\UARTTransmitter_ins.state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0185_));
 sky130_fd_sc_hd__a31o_1 _0569_ (.A1(net25),
    .A2(net59),
    .A3(_0181_),
    .B1(_0185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0005_));
 sky130_fd_sc_hd__a31o_1 _0570_ (.A1(\UARTTransmitter_ins.state[3] ),
    .A2(_0164_),
    .A3(_0165_),
    .B1(\UARTTransmitter_ins.state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0186_));
 sky130_fd_sc_hd__a21bo_1 _0571_ (.A1(net4),
    .A2(_0186_),
    .B1_N(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0004_));
 sky130_fd_sc_hd__nand4_4 _0572_ (.A(\UARTReceiver_ins.sampleCount[3] ),
    .B(\UARTReceiver_ins.sampleCount[2] ),
    .C(\UARTReceiver_ins.sampleCount[1] ),
    .D(\UARTReceiver_ins.sampleCount[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0187_));
 sky130_fd_sc_hd__o211a_1 _0573_ (.A1(_0152_),
    .A2(_0187_),
    .B1(net8),
    .C1(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0188_));
 sky130_fd_sc_hd__a31o_1 _0574_ (.A1(net19),
    .A2(net10),
    .A3(_0157_),
    .B1(_0188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0003_));
 sky130_fd_sc_hd__nor2_1 _0575_ (.A(_0148_),
    .B(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0189_));
 sky130_fd_sc_hd__nand2_1 _0576_ (.A(\UARTReceiver_ins.state[3] ),
    .B(_0143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0190_));
 sky130_fd_sc_hd__or4b_1 _0577_ (.A(\UARTReceiver_ins.sampleCount[2] ),
    .B(_0147_),
    .C(_0145_),
    .D_N(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0191_));
 sky130_fd_sc_hd__o21ai_1 _0578_ (.A1(_0142_),
    .A2(_0190_),
    .B1(_0191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0192_));
 sky130_fd_sc_hd__o21a_1 _0579_ (.A1(\UARTReceiver_ins.state[0] ),
    .A2(_0192_),
    .B1(_0155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0193_));
 sky130_fd_sc_hd__nor2_1 _0580_ (.A(_0147_),
    .B(_0155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0194_));
 sky130_fd_sc_hd__o31a_1 _0581_ (.A1(_0189_),
    .A2(_0193_),
    .A3(_0194_),
    .B1(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0002_));
 sky130_fd_sc_hd__and4bb_4 _0582_ (.A_N(\SRAMController_ins.cur_state[0] ),
    .B_N(\SRAMController_ins.cur_state[2] ),
    .C(\SRAMController_ins.cur_state[3] ),
    .D(\SRAMController_ins.cur_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0195_));
 sky130_fd_sc_hd__buf_2 _0583_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0196_));
 sky130_fd_sc_hd__and2_1 _0584_ (.A(\SRAMController_ins.data_tmp[0] ),
    .B(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0197_));
 sky130_fd_sc_hd__buf_1 _0585_ (.A(_0197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[0] ));
 sky130_fd_sc_hd__and2_1 _0586_ (.A(\SRAMController_ins.data_tmp[1] ),
    .B(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0198_));
 sky130_fd_sc_hd__buf_1 _0587_ (.A(_0198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[1] ));
 sky130_fd_sc_hd__and2_1 _0588_ (.A(\SRAMController_ins.data_tmp[2] ),
    .B(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0199_));
 sky130_fd_sc_hd__buf_1 _0589_ (.A(_0199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[2] ));
 sky130_fd_sc_hd__and2_1 _0590_ (.A(\SRAMController_ins.data_tmp[3] ),
    .B(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0200_));
 sky130_fd_sc_hd__buf_1 _0591_ (.A(_0200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[3] ));
 sky130_fd_sc_hd__and2_1 _0592_ (.A(\SRAMController_ins.data_tmp[4] ),
    .B(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0201_));
 sky130_fd_sc_hd__buf_1 _0593_ (.A(_0201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[4] ));
 sky130_fd_sc_hd__clkbuf_2 _0594_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0202_));
 sky130_fd_sc_hd__and2_1 _0595_ (.A(\SRAMController_ins.data_tmp[5] ),
    .B(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0203_));
 sky130_fd_sc_hd__buf_1 _0596_ (.A(_0203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[5] ));
 sky130_fd_sc_hd__and2_1 _0597_ (.A(\SRAMController_ins.data_tmp[6] ),
    .B(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0204_));
 sky130_fd_sc_hd__buf_1 _0598_ (.A(_0204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[6] ));
 sky130_fd_sc_hd__and2_1 _0599_ (.A(\SRAMController_ins.data_tmp[7] ),
    .B(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0205_));
 sky130_fd_sc_hd__buf_1 _0600_ (.A(_0205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[7] ));
 sky130_fd_sc_hd__and2_1 _0601_ (.A(\SRAMController_ins.data_tmp[8] ),
    .B(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0206_));
 sky130_fd_sc_hd__buf_1 _0602_ (.A(_0206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[8] ));
 sky130_fd_sc_hd__and2_1 _0603_ (.A(\SRAMController_ins.data_tmp[9] ),
    .B(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0207_));
 sky130_fd_sc_hd__buf_1 _0604_ (.A(_0207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[9] ));
 sky130_fd_sc_hd__and2_1 _0605_ (.A(\SRAMController_ins.data_tmp[10] ),
    .B(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0208_));
 sky130_fd_sc_hd__buf_1 _0606_ (.A(_0208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[10] ));
 sky130_fd_sc_hd__and2_1 _0607_ (.A(\SRAMController_ins.data_tmp[11] ),
    .B(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0209_));
 sky130_fd_sc_hd__buf_1 _0608_ (.A(_0209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[11] ));
 sky130_fd_sc_hd__and2_1 _0609_ (.A(\SRAMController_ins.data_tmp[12] ),
    .B(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0210_));
 sky130_fd_sc_hd__buf_1 _0610_ (.A(_0210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[12] ));
 sky130_fd_sc_hd__and2_1 _0611_ (.A(\SRAMController_ins.data_tmp[13] ),
    .B(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0211_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0612_ (.A(_0211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[13] ));
 sky130_fd_sc_hd__and2_1 _0613_ (.A(\SRAMController_ins.data_tmp[14] ),
    .B(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0212_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0614_ (.A(_0212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[14] ));
 sky130_fd_sc_hd__clkbuf_2 _0615_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0213_));
 sky130_fd_sc_hd__and2_1 _0616_ (.A(\SRAMController_ins.data_tmp[15] ),
    .B(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0214_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0617_ (.A(_0214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[15] ));
 sky130_fd_sc_hd__and2_1 _0618_ (.A(\SRAMController_ins.data_tmp[16] ),
    .B(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0215_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0619_ (.A(_0215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[16] ));
 sky130_fd_sc_hd__and2_1 _0620_ (.A(\SRAMController_ins.data_tmp[17] ),
    .B(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0216_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0621_ (.A(_0216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[17] ));
 sky130_fd_sc_hd__and2_1 _0622_ (.A(\SRAMController_ins.data_tmp[18] ),
    .B(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0217_));
 sky130_fd_sc_hd__clkbuf_2 _0623_ (.A(_0217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[18] ));
 sky130_fd_sc_hd__and2_1 _0624_ (.A(\SRAMController_ins.data_tmp[19] ),
    .B(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0218_));
 sky130_fd_sc_hd__clkbuf_2 _0625_ (.A(_0218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[19] ));
 sky130_fd_sc_hd__and2_1 _0626_ (.A(\SRAMController_ins.data_tmp[20] ),
    .B(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0219_));
 sky130_fd_sc_hd__clkbuf_2 _0627_ (.A(_0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[20] ));
 sky130_fd_sc_hd__and2_1 _0628_ (.A(\SRAMController_ins.data_tmp[21] ),
    .B(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_2 _0629_ (.A(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[21] ));
 sky130_fd_sc_hd__and2_1 _0630_ (.A(\SRAMController_ins.data_tmp[22] ),
    .B(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0221_));
 sky130_fd_sc_hd__clkbuf_2 _0631_ (.A(_0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[22] ));
 sky130_fd_sc_hd__and2_1 _0632_ (.A(\SRAMController_ins.data_tmp[23] ),
    .B(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_2 _0633_ (.A(_0222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[23] ));
 sky130_fd_sc_hd__and2_1 _0634_ (.A(\SRAMController_ins.data_tmp[24] ),
    .B(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0223_));
 sky130_fd_sc_hd__clkbuf_2 _0635_ (.A(_0223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[24] ));
 sky130_fd_sc_hd__and2_1 _0636_ (.A(\SRAMController_ins.data_tmp[25] ),
    .B(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0224_));
 sky130_fd_sc_hd__clkbuf_2 _0637_ (.A(_0224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[25] ));
 sky130_fd_sc_hd__and2_1 _0638_ (.A(\SRAMController_ins.data_tmp[26] ),
    .B(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0225_));
 sky130_fd_sc_hd__clkbuf_2 _0639_ (.A(_0225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[26] ));
 sky130_fd_sc_hd__and2_1 _0640_ (.A(\SRAMController_ins.data_tmp[27] ),
    .B(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_2 _0641_ (.A(_0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[27] ));
 sky130_fd_sc_hd__and2_1 _0642_ (.A(\SRAMController_ins.data_tmp[28] ),
    .B(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0227_));
 sky130_fd_sc_hd__clkbuf_2 _0643_ (.A(_0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[28] ));
 sky130_fd_sc_hd__and2_1 _0644_ (.A(\SRAMController_ins.data_tmp[29] ),
    .B(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0228_));
 sky130_fd_sc_hd__clkbuf_2 _0645_ (.A(_0228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[29] ));
 sky130_fd_sc_hd__and2_1 _0646_ (.A(\SRAMController_ins.data_tmp[30] ),
    .B(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0229_));
 sky130_fd_sc_hd__clkbuf_2 _0647_ (.A(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[30] ));
 sky130_fd_sc_hd__and2_1 _0648_ (.A(\SRAMController_ins.data_tmp[31] ),
    .B(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0230_));
 sky130_fd_sc_hd__buf_2 _0649_ (.A(_0230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.sram_data_in[31] ));
 sky130_fd_sc_hd__nor4_1 _0650_ (.A(\SRAMController_ins.cur_state[1] ),
    .B(\SRAMController_ins.cur_state[0] ),
    .C(\SRAMController_ins.cur_state[2] ),
    .D(\SRAMController_ins.cur_state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0231_));
 sky130_fd_sc_hd__and3_1 _0651_ (.A(\SRAMController_ins.rx_data_out[5] ),
    .B(\SRAMController_ins.rx_valid ),
    .C(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0232_));
 sky130_fd_sc_hd__clkbuf_4 _0652_ (.A(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.we_n ));
 sky130_fd_sc_hd__and2b_1 _0653_ (.A_N(net11),
    .B(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0233_));
 sky130_fd_sc_hd__or3b_1 _0654_ (.A(\SRAMController_ins.cur_state[1] ),
    .B(\SRAMController_ins.cur_state[2] ),
    .C_N(\SRAMController_ins.cur_state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0234_));
 sky130_fd_sc_hd__nand3b_1 _0655_ (.A_N(\SRAMController_ins.cur_state[3] ),
    .B(\SRAMController_ins.cur_state[2] ),
    .C(\SRAMController_ins.cur_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0235_));
 sky130_fd_sc_hd__nand2_1 _0656_ (.A(_0234_),
    .B(_0235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0236_));
 sky130_fd_sc_hd__nand2_1 _0657_ (.A(\SRAMController_ins.rx_valid ),
    .B(\SRAMController_ins.cur_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0237_));
 sky130_fd_sc_hd__or2_1 _0658_ (.A(\SRAMController_ins.rx_valid ),
    .B(\SRAMController_ins.cur_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0238_));
 sky130_fd_sc_hd__buf_6 _0659_ (.A(_0169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0239_));
 sky130_fd_sc_hd__and2b_1 _0660_ (.A_N(net11),
    .B(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0240_));
 sky130_fd_sc_hd__a31o_1 _0661_ (.A1(_0236_),
    .A2(_0237_),
    .A3(_0238_),
    .B1(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0241_));
 sky130_fd_sc_hd__nor2_1 _0662_ (.A(\SRAMController_ins.cur_state[0] ),
    .B(_0176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0242_));
 sky130_fd_sc_hd__or4_1 _0663_ (.A(\SRAMController_ins.we_n ),
    .B(_0233_),
    .C(_0241_),
    .D(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0243_));
 sky130_fd_sc_hd__clkbuf_1 _0664_ (.A(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.nxt_state[0] ));
 sky130_fd_sc_hd__inv_2 _0665_ (.A(\SRAMController_ins.cur_state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0244_));
 sky130_fd_sc_hd__and3b_2 _0666_ (.A_N(\SRAMController_ins.rx_data_out[5] ),
    .B(\SRAMController_ins.rx_valid ),
    .C(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0245_));
 sky130_fd_sc_hd__a41o_1 _0667_ (.A1(\SRAMController_ins.cur_state[1] ),
    .A2(\SRAMController_ins.cur_state[2] ),
    .A3(_0244_),
    .A4(_0237_),
    .B1(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0246_));
 sky130_fd_sc_hd__o21bai_1 _0668_ (.A1(_0234_),
    .A2(_0237_),
    .B1_N(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0247_));
 sky130_fd_sc_hd__or4b_1 _0669_ (.A(\SRAMController_ins.cur_state[1] ),
    .B(\SRAMController_ins.cur_state[2] ),
    .C(\SRAMController_ins.cur_state[3] ),
    .D_N(\SRAMController_ins.cur_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0248_));
 sky130_fd_sc_hd__buf_4 _0670_ (.A(_0248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0249_));
 sky130_fd_sc_hd__or4b_1 _0671_ (.A(_0240_),
    .B(_0246_),
    .C(_0247_),
    .D_N(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_1 _0672_ (.A(_0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.nxt_state[1] ));
 sky130_fd_sc_hd__a2111o_1 _0673_ (.A1(net11),
    .A2(_0239_),
    .B1(_0233_),
    .C1(_0246_),
    .D1(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.nxt_state[2] ));
 sky130_fd_sc_hd__o21ai_1 _0674_ (.A1(_0235_),
    .A2(_0237_),
    .B1(_0234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(\SRAMController_ins.nxt_state[3] ));
 sky130_fd_sc_hd__a22o_1 _0675_ (.A1(\SRAMController_ins.addr_tmp[0] ),
    .A2(_0196_),
    .B1(\SRAMController_ins.we_n ),
    .B2(\SRAMController_ins.rx_data_out[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.addr[0] ));
 sky130_fd_sc_hd__a22o_1 _0676_ (.A1(\SRAMController_ins.addr_tmp[1] ),
    .A2(_0196_),
    .B1(\SRAMController_ins.we_n ),
    .B2(\SRAMController_ins.rx_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.addr[1] ));
 sky130_fd_sc_hd__a22o_1 _0677_ (.A1(\SRAMController_ins.addr_tmp[2] ),
    .A2(_0196_),
    .B1(\SRAMController_ins.we_n ),
    .B2(\SRAMController_ins.rx_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.addr[2] ));
 sky130_fd_sc_hd__a22o_1 _0678_ (.A1(\SRAMController_ins.addr_tmp[3] ),
    .A2(_0196_),
    .B1(\SRAMController_ins.we_n ),
    .B2(\SRAMController_ins.rx_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(\SRAMController_ins.addr[3] ));
 sky130_fd_sc_hd__nor2_1 _0679_ (.A(_0196_),
    .B(\SRAMController_ins.we_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(\SRAMController_ins.csb_n ));
 sky130_fd_sc_hd__nor2_1 _0680_ (.A(net8),
    .B(\UARTReceiver_ins.state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0251_));
 sky130_fd_sc_hd__nand2_1 _0681_ (.A(_0147_),
    .B(_0251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0252_));
 sky130_fd_sc_hd__nand2_1 _0682_ (.A(_0148_),
    .B(_0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0253_));
 sky130_fd_sc_hd__o31ai_2 _0683_ (.A1(\SRAMController_ins.rx_valid ),
    .A2(_0142_),
    .A3(_0187_),
    .B1(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0254_));
 sky130_fd_sc_hd__a31o_1 _0684_ (.A1(_0148_),
    .A2(_0254_),
    .A3(_0252_),
    .B1(\UARTReceiver_ins.out_latched ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0255_));
 sky130_fd_sc_hd__o211a_1 _0685_ (.A1(net8),
    .A2(_0253_),
    .B1(_0255_),
    .C1(_0160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0008_));
 sky130_fd_sc_hd__a21oi_2 _0686_ (.A1(net10),
    .A2(_0187_),
    .B1(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0256_));
 sky130_fd_sc_hd__o2111ai_4 _0687_ (.A1(\UARTReceiver_ins.rxCounter[6] ),
    .A2(_0140_),
    .B1(_0148_),
    .C1(_0256_),
    .D1(\UARTReceiver_ins.rxCounter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0257_));
 sky130_fd_sc_hd__and2_1 _0688_ (.A(\UARTReceiver_ins.data[0] ),
    .B(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0258_));
 sky130_fd_sc_hd__o2111a_2 _0689_ (.A1(\UARTReceiver_ins.rxCounter[6] ),
    .A2(_0140_),
    .B1(_0148_),
    .C1(_0256_),
    .D1(\UARTReceiver_ins.rxCounter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0259_));
 sky130_fd_sc_hd__a21o_1 _0690_ (.A1(\UARTReceiver_ins.inputReg[1] ),
    .A2(\UARTReceiver_ins.inputReg[0] ),
    .B1(\UARTReceiver_ins.inputReg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0260_));
 sky130_fd_sc_hd__o21a_2 _0691_ (.A1(\UARTReceiver_ins.inputReg[1] ),
    .A2(\UARTReceiver_ins.inputReg[0] ),
    .B1(_0260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0261_));
 sky130_fd_sc_hd__or3_1 _0692_ (.A(\UARTReceiver_ins.bitIndex[2] ),
    .B(\UARTReceiver_ins.bitIndex[1] ),
    .C(\UARTReceiver_ins.bitIndex[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _0693_ (.A0(_0261_),
    .A1(\UARTReceiver_ins.data[0] ),
    .S(_0262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0263_));
 sky130_fd_sc_hd__and3_1 _0694_ (.A(net9),
    .B(_0259_),
    .C(_0263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0264_));
 sky130_fd_sc_hd__o21a_1 _0695_ (.A1(_0258_),
    .A2(_0264_),
    .B1(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0009_));
 sky130_fd_sc_hd__and2_1 _0696_ (.A(\UARTReceiver_ins.data[1] ),
    .B(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0265_));
 sky130_fd_sc_hd__inv_2 _0697_ (.A(\UARTReceiver_ins.bitIndex[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0266_));
 sky130_fd_sc_hd__or3_1 _0698_ (.A(\UARTReceiver_ins.bitIndex[2] ),
    .B(\UARTReceiver_ins.bitIndex[1] ),
    .C(_0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _0699_ (.A0(_0261_),
    .A1(\UARTReceiver_ins.data[1] ),
    .S(_0267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0268_));
 sky130_fd_sc_hd__and3_1 _0700_ (.A(net9),
    .B(_0259_),
    .C(_0268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0269_));
 sky130_fd_sc_hd__o21a_1 _0701_ (.A1(_0265_),
    .A2(_0269_),
    .B1(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0010_));
 sky130_fd_sc_hd__and2_1 _0702_ (.A(\UARTReceiver_ins.data[2] ),
    .B(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0270_));
 sky130_fd_sc_hd__or3b_1 _0703_ (.A(\UARTReceiver_ins.bitIndex[2] ),
    .B(\UARTReceiver_ins.bitIndex[0] ),
    .C_N(\UARTReceiver_ins.bitIndex[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _0704_ (.A0(_0261_),
    .A1(\UARTReceiver_ins.data[2] ),
    .S(_0271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0272_));
 sky130_fd_sc_hd__and3_1 _0705_ (.A(net9),
    .B(_0259_),
    .C(_0272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0273_));
 sky130_fd_sc_hd__o21a_1 _0706_ (.A1(_0270_),
    .A2(_0273_),
    .B1(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0011_));
 sky130_fd_sc_hd__and2_1 _0707_ (.A(\UARTReceiver_ins.data[3] ),
    .B(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0274_));
 sky130_fd_sc_hd__and2_1 _0708_ (.A(\UARTReceiver_ins.bitIndex[1] ),
    .B(\UARTReceiver_ins.bitIndex[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0275_));
 sky130_fd_sc_hd__and2b_1 _0709_ (.A_N(\UARTReceiver_ins.bitIndex[2] ),
    .B(_0275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _0710_ (.A0(\UARTReceiver_ins.data[3] ),
    .A1(_0261_),
    .S(_0276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0277_));
 sky130_fd_sc_hd__and3_1 _0711_ (.A(net9),
    .B(_0259_),
    .C(_0277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0278_));
 sky130_fd_sc_hd__o21a_1 _0712_ (.A1(_0274_),
    .A2(_0278_),
    .B1(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0012_));
 sky130_fd_sc_hd__and2_1 _0713_ (.A(\UARTReceiver_ins.data[4] ),
    .B(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0279_));
 sky130_fd_sc_hd__nor2_1 _0714_ (.A(\UARTReceiver_ins.bitIndex[1] ),
    .B(\UARTReceiver_ins.bitIndex[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0280_));
 sky130_fd_sc_hd__nand2_1 _0715_ (.A(\UARTReceiver_ins.bitIndex[2] ),
    .B(_0280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0281_));
 sky130_fd_sc_hd__mux2_1 _0716_ (.A0(_0261_),
    .A1(\UARTReceiver_ins.data[4] ),
    .S(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0282_));
 sky130_fd_sc_hd__and3_1 _0717_ (.A(net9),
    .B(_0259_),
    .C(_0282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0283_));
 sky130_fd_sc_hd__o21a_1 _0718_ (.A1(_0279_),
    .A2(_0283_),
    .B1(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0013_));
 sky130_fd_sc_hd__and2_1 _0719_ (.A(\UARTReceiver_ins.data[5] ),
    .B(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0284_));
 sky130_fd_sc_hd__and3b_1 _0720_ (.A_N(\UARTReceiver_ins.bitIndex[1] ),
    .B(\UARTReceiver_ins.bitIndex[0] ),
    .C(\UARTReceiver_ins.bitIndex[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _0721_ (.A0(\UARTReceiver_ins.data[5] ),
    .A1(_0261_),
    .S(_0285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0286_));
 sky130_fd_sc_hd__and3_1 _0722_ (.A(net9),
    .B(_0259_),
    .C(_0286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0287_));
 sky130_fd_sc_hd__o21a_1 _0723_ (.A1(_0284_),
    .A2(_0287_),
    .B1(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _0724_ (.A(\UARTReceiver_ins.data[6] ),
    .B(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0288_));
 sky130_fd_sc_hd__and3_1 _0725_ (.A(\UARTReceiver_ins.bitIndex[2] ),
    .B(\UARTReceiver_ins.bitIndex[1] ),
    .C(_0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _0726_ (.A0(\UARTReceiver_ins.data[6] ),
    .A1(_0261_),
    .S(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0290_));
 sky130_fd_sc_hd__and3_1 _0727_ (.A(net9),
    .B(_0259_),
    .C(_0290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0291_));
 sky130_fd_sc_hd__o21a_1 _0728_ (.A1(_0288_),
    .A2(_0291_),
    .B1(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0015_));
 sky130_fd_sc_hd__and2b_1 _0729_ (.A_N(_0156_),
    .B(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0292_));
 sky130_fd_sc_hd__o21a_1 _0730_ (.A1(_0257_),
    .A2(_0292_),
    .B1(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0293_));
 sky130_fd_sc_hd__and4_1 _0731_ (.A(net10),
    .B(_0156_),
    .C(_0259_),
    .D(_0261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0294_));
 sky130_fd_sc_hd__o21a_1 _0732_ (.A1(_0293_),
    .A2(_0294_),
    .B1(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0016_));
 sky130_fd_sc_hd__inv_2 _0733_ (.A(\UARTReceiver_ins.sampleCount[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0295_));
 sky130_fd_sc_hd__o21a_1 _0734_ (.A1(net10),
    .A2(_0252_),
    .B1(_0191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0296_));
 sky130_fd_sc_hd__nand2_1 _0735_ (.A(_0155_),
    .B(_0296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0297_));
 sky130_fd_sc_hd__nor2_1 _0736_ (.A(net8),
    .B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0298_));
 sky130_fd_sc_hd__nand2_1 _0737_ (.A(_0148_),
    .B(_0298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0299_));
 sky130_fd_sc_hd__a31o_1 _0738_ (.A1(_0155_),
    .A2(_0296_),
    .A3(_0299_),
    .B1(\UARTReceiver_ins.sampleCount[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0300_));
 sky130_fd_sc_hd__o211a_1 _0739_ (.A1(_0295_),
    .A2(_0297_),
    .B1(_0300_),
    .C1(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0017_));
 sky130_fd_sc_hd__a21boi_1 _0740_ (.A1(_0155_),
    .A2(_0296_),
    .B1_N(\UARTReceiver_ins.sampleCount[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0301_));
 sky130_fd_sc_hd__and2_1 _0741_ (.A(\UARTReceiver_ins.sampleCount[1] ),
    .B(\UARTReceiver_ins.sampleCount[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0302_));
 sky130_fd_sc_hd__nor2_1 _0742_ (.A(\UARTReceiver_ins.sampleCount[1] ),
    .B(\UARTReceiver_ins.sampleCount[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0303_));
 sky130_fd_sc_hd__nor2_1 _0743_ (.A(_0302_),
    .B(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0304_));
 sky130_fd_sc_hd__and4_1 _0744_ (.A(_0155_),
    .B(_0296_),
    .C(_0299_),
    .D(_0304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0305_));
 sky130_fd_sc_hd__o21a_1 _0745_ (.A1(_0301_),
    .A2(_0305_),
    .B1(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0018_));
 sky130_fd_sc_hd__a21boi_1 _0746_ (.A1(\UARTReceiver_ins.sampleCount[2] ),
    .A2(_0302_),
    .B1_N(_0299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0306_));
 sky130_fd_sc_hd__a31o_1 _0747_ (.A1(_0155_),
    .A2(_0302_),
    .A3(_0296_),
    .B1(\UARTReceiver_ins.sampleCount[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0307_));
 sky130_fd_sc_hd__o211a_1 _0748_ (.A1(_0297_),
    .A2(_0306_),
    .B1(_0307_),
    .C1(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0019_));
 sky130_fd_sc_hd__nor2_1 _0749_ (.A(_0143_),
    .B(_0298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0308_));
 sky130_fd_sc_hd__a31o_1 _0750_ (.A1(_0155_),
    .A2(_0302_),
    .A3(_0296_),
    .B1(\UARTReceiver_ins.sampleCount[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0309_));
 sky130_fd_sc_hd__o2111a_1 _0751_ (.A1(_0297_),
    .A2(_0308_),
    .B1(_0309_),
    .C1(net20),
    .D1(_0146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0020_));
 sky130_fd_sc_hd__o32a_1 _0752_ (.A1(\UARTReceiver_ins.state[0] ),
    .A2(net2),
    .A3(_0141_),
    .B1(_0153_),
    .B2(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0021_));
 sky130_fd_sc_hd__o32a_1 _0753_ (.A1(\UARTReceiver_ins.inputReg[0] ),
    .A2(\UARTReceiver_ins.state[0] ),
    .A3(_0141_),
    .B1(_0153_),
    .B2(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0022_));
 sky130_fd_sc_hd__o32a_1 _0754_ (.A1(\UARTReceiver_ins.inputReg[1] ),
    .A2(\UARTReceiver_ins.state[0] ),
    .A3(_0141_),
    .B1(_0153_),
    .B2(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0023_));
 sky130_fd_sc_hd__o211a_1 _0755_ (.A1(\UARTReceiver_ins.rxCounter[6] ),
    .A2(_0140_),
    .B1(_0148_),
    .C1(\UARTReceiver_ins.rxCounter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0310_));
 sky130_fd_sc_hd__nand2_1 _0756_ (.A(net10),
    .B(_0187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0311_));
 sky130_fd_sc_hd__o31a_1 _0757_ (.A1(\UARTReceiver_ins.state[0] ),
    .A2(\UARTReceiver_ins.state[2] ),
    .A3(net10),
    .B1(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0312_));
 sky130_fd_sc_hd__nand2_1 _0758_ (.A(_0310_),
    .B(_0312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0313_));
 sky130_fd_sc_hd__a31o_1 _0759_ (.A1(net9),
    .A2(_0310_),
    .A3(_0311_),
    .B1(\UARTReceiver_ins.bitIndex[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0314_));
 sky130_fd_sc_hd__o211a_1 _0760_ (.A1(_0266_),
    .A2(_0313_),
    .B1(_0314_),
    .C1(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0024_));
 sky130_fd_sc_hd__a21boi_1 _0761_ (.A1(_0310_),
    .A2(_0312_),
    .B1_N(\UARTReceiver_ins.bitIndex[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0315_));
 sky130_fd_sc_hd__nor2_1 _0762_ (.A(_0275_),
    .B(_0280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0316_));
 sky130_fd_sc_hd__and4_1 _0763_ (.A(net9),
    .B(_0310_),
    .C(_0311_),
    .D(_0316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0317_));
 sky130_fd_sc_hd__o21a_1 _0764_ (.A1(_0315_),
    .A2(_0317_),
    .B1(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0025_));
 sky130_fd_sc_hd__a41o_1 _0765_ (.A1(\UARTReceiver_ins.bitIndex[1] ),
    .A2(\UARTReceiver_ins.bitIndex[0] ),
    .A3(_0310_),
    .A4(_0312_),
    .B1(\UARTReceiver_ins.bitIndex[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0318_));
 sky130_fd_sc_hd__o211a_1 _0766_ (.A1(_0292_),
    .A2(_0313_),
    .B1(_0318_),
    .C1(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _0767_ (.A0(\SRAMController_ins.addr_tmp[0] ),
    .A1(\SRAMController_ins.rx_data_out[0] ),
    .S(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_1 _0768_ (.A(_0319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _0769_ (.A0(\SRAMController_ins.addr_tmp[1] ),
    .A1(\SRAMController_ins.rx_data_out[1] ),
    .S(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_1 _0770_ (.A(_0320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _0771_ (.A0(\SRAMController_ins.addr_tmp[2] ),
    .A1(\SRAMController_ins.rx_data_out[2] ),
    .S(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _0772_ (.A(_0321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _0773_ (.A0(\SRAMController_ins.addr_tmp[3] ),
    .A1(\SRAMController_ins.rx_data_out[3] ),
    .S(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0322_));
 sky130_fd_sc_hd__clkbuf_1 _0774_ (.A(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0030_));
 sky130_fd_sc_hd__nand2_1 _0775_ (.A(net8),
    .B(_0187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0323_));
 sky130_fd_sc_hd__or2b_1 _0776_ (.A(\SRAMController_ins.rx_valid ),
    .B_N(\UARTReceiver_ins.state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0324_));
 sky130_fd_sc_hd__and4b_1 _0777_ (.A_N(_0144_),
    .B(_0148_),
    .C(_0252_),
    .D(_0324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0325_));
 sky130_fd_sc_hd__a31o_1 _0778_ (.A1(_0154_),
    .A2(_0323_),
    .A3(_0325_),
    .B1(\UARTReceiver_ins.overrun ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0326_));
 sky130_fd_sc_hd__or3b_1 _0779_ (.A(net8),
    .B(_0152_),
    .C_N(_0325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0327_));
 sky130_fd_sc_hd__and3_1 _0780_ (.A(net17),
    .B(_0326_),
    .C(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_1 _0781_ (.A(_0328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0031_));
 sky130_fd_sc_hd__o21a_1 _0782_ (.A1(_0148_),
    .A2(_0149_),
    .B1(_0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0329_));
 sky130_fd_sc_hd__and4bb_1 _0783_ (.A_N(_0152_),
    .B_N(_0192_),
    .C(_0323_),
    .D(_0329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0330_));
 sky130_fd_sc_hd__o211a_1 _0784_ (.A1(net73),
    .A2(_0330_),
    .B1(_0327_),
    .C1(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0032_));
 sky130_fd_sc_hd__o21a_1 _0785_ (.A1(\UARTReceiver_ins.state[0] ),
    .A2(_0152_),
    .B1(\UARTReceiver_ins.out_latched ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0331_));
 sky130_fd_sc_hd__nor2_1 _0786_ (.A(net5),
    .B(_0236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0332_));
 sky130_fd_sc_hd__o211a_1 _0787_ (.A1(\UARTReceiver_ins.out_latched ),
    .A2(_0332_),
    .B1(_0152_),
    .C1(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0333_));
 sky130_fd_sc_hd__nor2_1 _0788_ (.A(\UARTReceiver_ins.state[0] ),
    .B(_0141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0334_));
 sky130_fd_sc_hd__o22a_1 _0789_ (.A1(net84),
    .A2(_0331_),
    .B1(_0333_),
    .B2(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0033_));
 sky130_fd_sc_hd__inv_2 _0790_ (.A(_0254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0335_));
 sky130_fd_sc_hd__o31a_2 _0791_ (.A1(_0152_),
    .A2(_0335_),
    .A3(_0251_),
    .B1(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0336_));
 sky130_fd_sc_hd__and4_1 _0792_ (.A(net8),
    .B(net19),
    .C(_0154_),
    .D(_0254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_2 _0793_ (.A(_0337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0338_));
 sky130_fd_sc_hd__a22o_1 _0794_ (.A1(\SRAMController_ins.rx_data_out[0] ),
    .A2(_0336_),
    .B1(_0338_),
    .B2(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0034_));
 sky130_fd_sc_hd__a22o_1 _0795_ (.A1(\SRAMController_ins.rx_data_out[1] ),
    .A2(_0336_),
    .B1(_0338_),
    .B2(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0035_));
 sky130_fd_sc_hd__a22o_1 _0796_ (.A1(\SRAMController_ins.rx_data_out[2] ),
    .A2(_0336_),
    .B1(_0338_),
    .B2(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0036_));
 sky130_fd_sc_hd__a22o_1 _0797_ (.A1(\SRAMController_ins.rx_data_out[3] ),
    .A2(_0336_),
    .B1(_0338_),
    .B2(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0037_));
 sky130_fd_sc_hd__a22o_1 _0798_ (.A1(\SRAMController_ins.rx_data_out[4] ),
    .A2(_0336_),
    .B1(_0338_),
    .B2(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0038_));
 sky130_fd_sc_hd__a22o_1 _0799_ (.A1(\SRAMController_ins.rx_data_out[5] ),
    .A2(_0336_),
    .B1(_0338_),
    .B2(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0039_));
 sky130_fd_sc_hd__a22o_1 _0800_ (.A1(\SRAMController_ins.rx_data_out[6] ),
    .A2(_0336_),
    .B1(_0338_),
    .B2(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0040_));
 sky130_fd_sc_hd__a22o_1 _0801_ (.A1(\SRAMController_ins.rx_data_out[7] ),
    .A2(_0336_),
    .B1(_0338_),
    .B2(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0041_));
 sky130_fd_sc_hd__nand2_1 _0802_ (.A(\UARTTransmitter_ins.txCounter[0] ),
    .B(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0339_));
 sky130_fd_sc_hd__o211a_1 _0803_ (.A1(\UARTTransmitter_ins.txCounter[0] ),
    .A2(_0172_),
    .B1(_0339_),
    .C1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0042_));
 sky130_fd_sc_hd__xnor2_1 _0804_ (.A(\UARTTransmitter_ins.txCounter[1] ),
    .B(_0339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0340_));
 sky130_fd_sc_hd__and2_1 _0805_ (.A(_0182_),
    .B(_0340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0341_));
 sky130_fd_sc_hd__clkbuf_1 _0806_ (.A(_0341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0043_));
 sky130_fd_sc_hd__and3_1 _0807_ (.A(\UARTTransmitter_ins.txCounter[2] ),
    .B(\UARTTransmitter_ins.txCounter[1] ),
    .C(\UARTTransmitter_ins.txCounter[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0342_));
 sky130_fd_sc_hd__inv_2 _0808_ (.A(_0342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0343_));
 sky130_fd_sc_hd__a32o_1 _0809_ (.A1(_0161_),
    .A2(_0172_),
    .A3(_0343_),
    .B1(_0171_),
    .B2(\UARTTransmitter_ins.txCounter[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0344_));
 sky130_fd_sc_hd__and2_1 _0810_ (.A(net26),
    .B(_0344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_1 _0811_ (.A(_0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0044_));
 sky130_fd_sc_hd__and4_2 _0812_ (.A(\UARTTransmitter_ins.txCounter[3] ),
    .B(\UARTTransmitter_ins.txCounter[2] ),
    .C(\UARTTransmitter_ins.txCounter[1] ),
    .D(\UARTTransmitter_ins.txCounter[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0346_));
 sky130_fd_sc_hd__inv_2 _0813_ (.A(_0346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0347_));
 sky130_fd_sc_hd__a22o_1 _0814_ (.A1(\UARTTransmitter_ins.txCounter[3] ),
    .A2(_0171_),
    .B1(_0172_),
    .B2(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0348_));
 sky130_fd_sc_hd__o211a_1 _0815_ (.A1(\UARTTransmitter_ins.txCounter[3] ),
    .A2(_0342_),
    .B1(_0348_),
    .C1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0045_));
 sky130_fd_sc_hd__nand2_1 _0816_ (.A(\UARTTransmitter_ins.txCounter[4] ),
    .B(_0346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0349_));
 sky130_fd_sc_hd__a22o_1 _0817_ (.A1(\UARTTransmitter_ins.txCounter[4] ),
    .A2(_0171_),
    .B1(_0172_),
    .B2(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0350_));
 sky130_fd_sc_hd__o211a_1 _0818_ (.A1(\UARTTransmitter_ins.txCounter[4] ),
    .A2(_0346_),
    .B1(_0350_),
    .C1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0046_));
 sky130_fd_sc_hd__a21o_1 _0819_ (.A1(\UARTTransmitter_ins.txCounter[4] ),
    .A2(_0346_),
    .B1(\UARTTransmitter_ins.txCounter[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0351_));
 sky130_fd_sc_hd__and2_1 _0820_ (.A(_0163_),
    .B(_0346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0352_));
 sky130_fd_sc_hd__inv_2 _0821_ (.A(_0352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0353_));
 sky130_fd_sc_hd__a22o_1 _0822_ (.A1(\UARTTransmitter_ins.txCounter[5] ),
    .A2(_0171_),
    .B1(_0172_),
    .B2(_0353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0354_));
 sky130_fd_sc_hd__and3_1 _0823_ (.A(net26),
    .B(_0351_),
    .C(_0354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_1 _0824_ (.A(_0355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0047_));
 sky130_fd_sc_hd__nand2_1 _0825_ (.A(\UARTTransmitter_ins.txCounter[6] ),
    .B(_0352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0356_));
 sky130_fd_sc_hd__a22o_1 _0826_ (.A1(\UARTTransmitter_ins.txCounter[6] ),
    .A2(_0171_),
    .B1(_0172_),
    .B2(_0356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0357_));
 sky130_fd_sc_hd__o211a_1 _0827_ (.A1(\UARTTransmitter_ins.txCounter[6] ),
    .A2(_0352_),
    .B1(_0357_),
    .C1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0048_));
 sky130_fd_sc_hd__a31o_1 _0828_ (.A1(\UARTTransmitter_ins.txCounter[6] ),
    .A2(_0163_),
    .A3(_0346_),
    .B1(\UARTTransmitter_ins.txCounter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0358_));
 sky130_fd_sc_hd__and4_1 _0829_ (.A(\UARTTransmitter_ins.txCounter[7] ),
    .B(\UARTTransmitter_ins.txCounter[6] ),
    .C(_0163_),
    .D(_0346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0359_));
 sky130_fd_sc_hd__inv_2 _0830_ (.A(_0359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0360_));
 sky130_fd_sc_hd__a22o_1 _0831_ (.A1(\UARTTransmitter_ins.txCounter[7] ),
    .A2(_0171_),
    .B1(_0172_),
    .B2(_0360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0361_));
 sky130_fd_sc_hd__and3_1 _0832_ (.A(net26),
    .B(_0358_),
    .C(_0361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_1 _0833_ (.A(_0362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0049_));
 sky130_fd_sc_hd__and3_1 _0834_ (.A(\UARTTransmitter_ins.txCounter[8] ),
    .B(net3),
    .C(_0359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0363_));
 sky130_fd_sc_hd__a21o_1 _0835_ (.A1(_0172_),
    .A2(_0359_),
    .B1(\UARTTransmitter_ins.txCounter[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0364_));
 sky130_fd_sc_hd__and3b_1 _0836_ (.A_N(_0363_),
    .B(_0182_),
    .C(_0364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_1 _0837_ (.A(_0365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0050_));
 sky130_fd_sc_hd__or2_1 _0838_ (.A(\UARTTransmitter_ins.txCounter[9] ),
    .B(_0363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0366_));
 sky130_fd_sc_hd__nand2_1 _0839_ (.A(\UARTTransmitter_ins.txCounter[9] ),
    .B(_0363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0367_));
 sky130_fd_sc_hd__and3_1 _0840_ (.A(_0182_),
    .B(_0366_),
    .C(_0367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_1 _0841_ (.A(_0368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0051_));
 sky130_fd_sc_hd__a21o_1 _0842_ (.A1(\UARTTransmitter_ins.txCounter[9] ),
    .A2(_0363_),
    .B1(\UARTTransmitter_ins.txCounter[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0369_));
 sky130_fd_sc_hd__nand3_1 _0843_ (.A(\UARTTransmitter_ins.txCounter[10] ),
    .B(\UARTTransmitter_ins.txCounter[9] ),
    .C(_0363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0370_));
 sky130_fd_sc_hd__and3_1 _0844_ (.A(_0182_),
    .B(_0369_),
    .C(_0370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0371_));
 sky130_fd_sc_hd__clkbuf_1 _0845_ (.A(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0052_));
 sky130_fd_sc_hd__inv_2 _0846_ (.A(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0372_));
 sky130_fd_sc_hd__a21boi_1 _0847_ (.A1(_0372_),
    .A2(_0370_),
    .B1_N(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0053_));
 sky130_fd_sc_hd__a31o_1 _0848_ (.A1(\UARTTransmitter_ins.state[0] ),
    .A2(_0164_),
    .A3(_0165_),
    .B1(_0170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0373_));
 sky130_fd_sc_hd__buf_2 _0849_ (.A(_0373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0374_));
 sky130_fd_sc_hd__a22o_1 _0850_ (.A1(\SRAMController_ins.sram_tmp[0] ),
    .A2(_0173_),
    .B1(_0175_),
    .B2(\SRAMController_ins.sram_tmp[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0375_));
 sky130_fd_sc_hd__a221o_4 _0851_ (.A1(\SRAMController_ins.sram_tmp[16] ),
    .A2(_0174_),
    .B1(_0239_),
    .B2(\SRAMController_ins.sram_tmp[8] ),
    .C1(_0375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0376_));
 sky130_fd_sc_hd__a21bo_1 _0852_ (.A1(\SRAMController_ins.tx_ready ),
    .A2(_0376_),
    .B1_N(_0374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0377_));
 sky130_fd_sc_hd__o211a_1 _0853_ (.A1(net67),
    .A2(_0374_),
    .B1(_0377_),
    .C1(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0054_));
 sky130_fd_sc_hd__a22o_1 _0854_ (.A1(\SRAMController_ins.sram_tmp[25] ),
    .A2(_0175_),
    .B1(_0239_),
    .B2(\SRAMController_ins.sram_tmp[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0378_));
 sky130_fd_sc_hd__a221o_1 _0855_ (.A1(\SRAMController_ins.sram_tmp[1] ),
    .A2(_0173_),
    .B1(_0174_),
    .B2(\SRAMController_ins.sram_tmp[17] ),
    .C1(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0379_));
 sky130_fd_sc_hd__a21bo_1 _0856_ (.A1(net11),
    .A2(_0379_),
    .B1_N(_0374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0380_));
 sky130_fd_sc_hd__o211a_1 _0857_ (.A1(net68),
    .A2(_0374_),
    .B1(_0380_),
    .C1(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0055_));
 sky130_fd_sc_hd__a22o_1 _0858_ (.A1(\SRAMController_ins.sram_tmp[26] ),
    .A2(_0175_),
    .B1(_0239_),
    .B2(\SRAMController_ins.sram_tmp[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0381_));
 sky130_fd_sc_hd__a221o_4 _0859_ (.A1(\SRAMController_ins.sram_tmp[2] ),
    .A2(_0173_),
    .B1(_0174_),
    .B2(\SRAMController_ins.sram_tmp[18] ),
    .C1(_0381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0382_));
 sky130_fd_sc_hd__a21bo_1 _0860_ (.A1(\SRAMController_ins.tx_ready ),
    .A2(_0382_),
    .B1_N(_0374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0383_));
 sky130_fd_sc_hd__o211a_1 _0861_ (.A1(net71),
    .A2(_0374_),
    .B1(_0383_),
    .C1(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0056_));
 sky130_fd_sc_hd__inv_2 _0862_ (.A(\UARTTransmitter_ins.data[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0384_));
 sky130_fd_sc_hd__a22o_1 _0863_ (.A1(\SRAMController_ins.sram_tmp[27] ),
    .A2(_0175_),
    .B1(_0239_),
    .B2(\SRAMController_ins.sram_tmp[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0385_));
 sky130_fd_sc_hd__a221o_2 _0864_ (.A1(\SRAMController_ins.sram_tmp[3] ),
    .A2(_0173_),
    .B1(_0174_),
    .B2(\SRAMController_ins.sram_tmp[19] ),
    .C1(_0385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0386_));
 sky130_fd_sc_hd__a2bb2o_1 _0865_ (.A1_N(_0384_),
    .A2_N(_0373_),
    .B1(_0386_),
    .B2(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0387_));
 sky130_fd_sc_hd__and2_1 _0866_ (.A(net22),
    .B(_0387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0388_));
 sky130_fd_sc_hd__clkbuf_1 _0867_ (.A(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0057_));
 sky130_fd_sc_hd__inv_2 _0868_ (.A(\UARTTransmitter_ins.data[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0389_));
 sky130_fd_sc_hd__a22o_1 _0869_ (.A1(\SRAMController_ins.sram_tmp[28] ),
    .A2(_0175_),
    .B1(_0239_),
    .B2(\SRAMController_ins.sram_tmp[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0390_));
 sky130_fd_sc_hd__a221o_2 _0870_ (.A1(\SRAMController_ins.sram_tmp[4] ),
    .A2(_0173_),
    .B1(_0174_),
    .B2(\SRAMController_ins.sram_tmp[20] ),
    .C1(_0390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0391_));
 sky130_fd_sc_hd__a2bb2o_1 _0871_ (.A1_N(_0389_),
    .A2_N(_0373_),
    .B1(_0391_),
    .B2(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0392_));
 sky130_fd_sc_hd__and2_1 _0872_ (.A(net25),
    .B(_0392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _0873_ (.A(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0058_));
 sky130_fd_sc_hd__a22o_1 _0874_ (.A1(\SRAMController_ins.sram_tmp[29] ),
    .A2(_0175_),
    .B1(_0239_),
    .B2(\SRAMController_ins.sram_tmp[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0394_));
 sky130_fd_sc_hd__a221o_2 _0875_ (.A1(\SRAMController_ins.sram_tmp[5] ),
    .A2(_0173_),
    .B1(_0174_),
    .B2(\SRAMController_ins.sram_tmp[21] ),
    .C1(_0394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0395_));
 sky130_fd_sc_hd__a21bo_1 _0876_ (.A1(net11),
    .A2(_0395_),
    .B1_N(_0374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0396_));
 sky130_fd_sc_hd__o211a_1 _0877_ (.A1(net65),
    .A2(_0374_),
    .B1(_0396_),
    .C1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0059_));
 sky130_fd_sc_hd__a22o_1 _0878_ (.A1(\SRAMController_ins.sram_tmp[6] ),
    .A2(_0173_),
    .B1(_0175_),
    .B2(\SRAMController_ins.sram_tmp[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0397_));
 sky130_fd_sc_hd__a221o_1 _0879_ (.A1(\SRAMController_ins.sram_tmp[22] ),
    .A2(_0174_),
    .B1(_0239_),
    .B2(\SRAMController_ins.sram_tmp[14] ),
    .C1(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0398_));
 sky130_fd_sc_hd__inv_2 _0880_ (.A(\UARTTransmitter_ins.data[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0399_));
 sky130_fd_sc_hd__o2bb2a_1 _0881_ (.A1_N(\SRAMController_ins.tx_ready ),
    .A2_N(_0398_),
    .B1(_0373_),
    .B2(_0399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0400_));
 sky130_fd_sc_hd__and2b_1 _0882_ (.A_N(_0400_),
    .B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _0883_ (.A(_0401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0060_));
 sky130_fd_sc_hd__a22o_1 _0884_ (.A1(\SRAMController_ins.sram_tmp[31] ),
    .A2(_0175_),
    .B1(_0239_),
    .B2(\SRAMController_ins.sram_tmp[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0402_));
 sky130_fd_sc_hd__a221o_2 _0885_ (.A1(\SRAMController_ins.sram_tmp[7] ),
    .A2(_0173_),
    .B1(_0174_),
    .B2(\SRAMController_ins.sram_tmp[23] ),
    .C1(_0402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0403_));
 sky130_fd_sc_hd__a21bo_1 _0886_ (.A1(\SRAMController_ins.tx_ready ),
    .A2(_0403_),
    .B1_N(_0374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0404_));
 sky130_fd_sc_hd__o211a_1 _0887_ (.A1(net66),
    .A2(_0374_),
    .B1(_0404_),
    .C1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0061_));
 sky130_fd_sc_hd__nor2_1 _0888_ (.A(\UARTTransmitter_ins.state[0] ),
    .B(\UARTTransmitter_ins.state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0405_));
 sky130_fd_sc_hd__nand3b_1 _0889_ (.A_N(_0405_),
    .B(_0181_),
    .C(\UARTTransmitter_ins.bitIndex[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0406_));
 sky130_fd_sc_hd__o211a_1 _0890_ (.A1(\UARTTransmitter_ins.bitIndex[0] ),
    .A2(_0177_),
    .B1(_0406_),
    .C1(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0062_));
 sky130_fd_sc_hd__o31a_1 _0891_ (.A1(_0183_),
    .A2(_0171_),
    .A3(_0405_),
    .B1(\UARTTransmitter_ins.bitIndex[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0407_));
 sky130_fd_sc_hd__nand2_1 _0892_ (.A(\UARTTransmitter_ins.bitIndex[1] ),
    .B(\UARTTransmitter_ins.bitIndex[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0408_));
 sky130_fd_sc_hd__or2_1 _0893_ (.A(\UARTTransmitter_ins.bitIndex[1] ),
    .B(\UARTTransmitter_ins.bitIndex[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0409_));
 sky130_fd_sc_hd__and3_1 _0894_ (.A(_0177_),
    .B(_0408_),
    .C(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0410_));
 sky130_fd_sc_hd__o21a_1 _0895_ (.A1(_0407_),
    .A2(_0410_),
    .B1(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0063_));
 sky130_fd_sc_hd__o31a_1 _0896_ (.A1(_0183_),
    .A2(_0171_),
    .A3(_0405_),
    .B1(\UARTTransmitter_ins.bitIndex[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0411_));
 sky130_fd_sc_hd__a21o_1 _0897_ (.A1(\UARTTransmitter_ins.bitIndex[1] ),
    .A2(\UARTTransmitter_ins.bitIndex[0] ),
    .B1(\UARTTransmitter_ins.bitIndex[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0412_));
 sky130_fd_sc_hd__and3_1 _0898_ (.A(_0177_),
    .B(_0184_),
    .C(_0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0413_));
 sky130_fd_sc_hd__o21a_1 _0899_ (.A1(_0411_),
    .A2(_0413_),
    .B1(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0064_));
 sky130_fd_sc_hd__inv_2 _0900_ (.A(\UARTTransmitter_ins.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0414_));
 sky130_fd_sc_hd__nand2_1 _0901_ (.A(net24),
    .B(_0181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0415_));
 sky130_fd_sc_hd__mux4_1 _0902_ (.A0(\UARTTransmitter_ins.data[0] ),
    .A1(\UARTTransmitter_ins.data[1] ),
    .A2(\UARTTransmitter_ins.data[2] ),
    .A3(\UARTTransmitter_ins.data[3] ),
    .S0(\UARTTransmitter_ins.bitIndex[0] ),
    .S1(\UARTTransmitter_ins.bitIndex[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0416_));
 sky130_fd_sc_hd__mux4_1 _0903_ (.A0(\UARTTransmitter_ins.data[4] ),
    .A1(\UARTTransmitter_ins.data[5] ),
    .A2(\UARTTransmitter_ins.data[6] ),
    .A3(\UARTTransmitter_ins.data[7] ),
    .S0(\UARTTransmitter_ins.bitIndex[0] ),
    .S1(\UARTTransmitter_ins.bitIndex[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _0904_ (.A0(_0416_),
    .A1(_0417_),
    .S(\UARTTransmitter_ins.bitIndex[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0418_));
 sky130_fd_sc_hd__a211o_1 _0905_ (.A1(\UARTTransmitter_ins.state[1] ),
    .A2(_0418_),
    .B1(\UARTTransmitter_ins.state[3] ),
    .C1(\UARTTransmitter_ins.state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0419_));
 sky130_fd_sc_hd__o2bb2a_1 _0906_ (.A1_N(_0414_),
    .A2_N(_0182_),
    .B1(_0415_),
    .B2(_0419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0065_));
 sky130_fd_sc_hd__a31o_1 _0907_ (.A1(\UARTTransmitter_ins.state[0] ),
    .A2(_0164_),
    .A3(_0165_),
    .B1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0420_));
 sky130_fd_sc_hd__and3_1 _0908_ (.A(net24),
    .B(net4),
    .C(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_1 _0909_ (.A(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0066_));
 sky130_fd_sc_hd__nor2_1 _0910_ (.A(net60),
    .B(_0153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0067_));
 sky130_fd_sc_hd__and2_1 _0911_ (.A(net21),
    .B(_0152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0422_));
 sky130_fd_sc_hd__nand2_1 _0912_ (.A(\UARTReceiver_ins.rxCounter[0] ),
    .B(\UARTReceiver_ins.rxCounter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0423_));
 sky130_fd_sc_hd__and3_1 _0913_ (.A(_0139_),
    .B(_0422_),
    .C(_0423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_1 _0914_ (.A(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0068_));
 sky130_fd_sc_hd__and3_1 _0915_ (.A(\UARTReceiver_ins.rxCounter[0] ),
    .B(\UARTReceiver_ins.rxCounter[2] ),
    .C(\UARTReceiver_ins.rxCounter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0425_));
 sky130_fd_sc_hd__a21o_1 _0916_ (.A1(\UARTReceiver_ins.rxCounter[0] ),
    .A2(\UARTReceiver_ins.rxCounter[1] ),
    .B1(\UARTReceiver_ins.rxCounter[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0426_));
 sky130_fd_sc_hd__and3b_1 _0917_ (.A_N(_0425_),
    .B(_0426_),
    .C(_0422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_1 _0918_ (.A(_0427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0069_));
 sky130_fd_sc_hd__and2_1 _0919_ (.A(\UARTReceiver_ins.rxCounter[3] ),
    .B(_0425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0428_));
 sky130_fd_sc_hd__or2_1 _0920_ (.A(\UARTReceiver_ins.rxCounter[3] ),
    .B(_0425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0429_));
 sky130_fd_sc_hd__and3b_1 _0921_ (.A_N(_0428_),
    .B(_0429_),
    .C(_0422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _0922_ (.A(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0070_));
 sky130_fd_sc_hd__and3_1 _0923_ (.A(\UARTReceiver_ins.rxCounter[4] ),
    .B(\UARTReceiver_ins.rxCounter[3] ),
    .C(_0425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0431_));
 sky130_fd_sc_hd__or2_1 _0924_ (.A(\UARTReceiver_ins.rxCounter[4] ),
    .B(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0432_));
 sky130_fd_sc_hd__and3b_1 _0925_ (.A_N(_0431_),
    .B(_0432_),
    .C(_0422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_1 _0926_ (.A(_0433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0071_));
 sky130_fd_sc_hd__and3_1 _0927_ (.A(\UARTReceiver_ins.rxCounter[5] ),
    .B(\UARTReceiver_ins.rxCounter[4] ),
    .C(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0434_));
 sky130_fd_sc_hd__or2_1 _0928_ (.A(\UARTReceiver_ins.rxCounter[5] ),
    .B(_0431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0435_));
 sky130_fd_sc_hd__and3b_1 _0929_ (.A_N(_0434_),
    .B(_0435_),
    .C(_0422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _0930_ (.A(_0436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0072_));
 sky130_fd_sc_hd__nand2_1 _0931_ (.A(\UARTReceiver_ins.rxCounter[6] ),
    .B(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0437_));
 sky130_fd_sc_hd__or2_1 _0932_ (.A(\UARTReceiver_ins.rxCounter[6] ),
    .B(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0438_));
 sky130_fd_sc_hd__and3_1 _0933_ (.A(_0422_),
    .B(_0437_),
    .C(_0438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0439_));
 sky130_fd_sc_hd__clkbuf_1 _0934_ (.A(_0439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0073_));
 sky130_fd_sc_hd__inv_2 _0935_ (.A(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0440_));
 sky130_fd_sc_hd__a21oi_1 _0936_ (.A1(_0440_),
    .A2(_0437_),
    .B1(_0153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Y(_0074_));
 sky130_fd_sc_hd__clkbuf_8 _0937_ (.A(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _0938_ (.A0(\SRAMController_ins.sram_data_out[0] ),
    .A1(\SRAMController_ins.sram_tmp[0] ),
    .S(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _0939_ (.A(_0442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _0940_ (.A0(\SRAMController_ins.sram_data_out[1] ),
    .A1(\SRAMController_ins.sram_tmp[1] ),
    .S(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_1 _0941_ (.A(_0443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _0942_ (.A0(\SRAMController_ins.sram_data_out[2] ),
    .A1(\SRAMController_ins.sram_tmp[2] ),
    .S(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_1 _0943_ (.A(_0444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _0944_ (.A0(\SRAMController_ins.sram_data_out[3] ),
    .A1(\SRAMController_ins.sram_tmp[3] ),
    .S(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_1 _0945_ (.A(_0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0946_ (.A0(\SRAMController_ins.sram_data_out[4] ),
    .A1(\SRAMController_ins.sram_tmp[4] ),
    .S(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _0947_ (.A(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _0948_ (.A0(\SRAMController_ins.sram_data_out[5] ),
    .A1(\SRAMController_ins.sram_tmp[5] ),
    .S(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _0949_ (.A(_0447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _0950_ (.A0(\SRAMController_ins.sram_data_out[6] ),
    .A1(\SRAMController_ins.sram_tmp[6] ),
    .S(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _0951_ (.A(_0448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _0952_ (.A0(\SRAMController_ins.sram_data_out[7] ),
    .A1(\SRAMController_ins.sram_tmp[7] ),
    .S(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _0953_ (.A(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _0954_ (.A0(\SRAMController_ins.sram_data_out[8] ),
    .A1(\SRAMController_ins.sram_tmp[8] ),
    .S(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_1 _0955_ (.A(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _0956_ (.A0(\SRAMController_ins.sram_data_out[9] ),
    .A1(\SRAMController_ins.sram_tmp[9] ),
    .S(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_1 _0957_ (.A(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0084_));
 sky130_fd_sc_hd__buf_6 _0958_ (.A(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _0959_ (.A0(\SRAMController_ins.sram_data_out[10] ),
    .A1(\SRAMController_ins.sram_tmp[10] ),
    .S(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0453_));
 sky130_fd_sc_hd__clkbuf_1 _0960_ (.A(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _0961_ (.A0(\SRAMController_ins.sram_data_out[11] ),
    .A1(\SRAMController_ins.sram_tmp[11] ),
    .S(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_1 _0962_ (.A(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _0963_ (.A0(\SRAMController_ins.sram_data_out[12] ),
    .A1(\SRAMController_ins.sram_tmp[12] ),
    .S(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_1 _0964_ (.A(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _0965_ (.A0(\SRAMController_ins.sram_data_out[13] ),
    .A1(\SRAMController_ins.sram_tmp[13] ),
    .S(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_1 _0966_ (.A(_0456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _0967_ (.A0(\SRAMController_ins.sram_data_out[14] ),
    .A1(\SRAMController_ins.sram_tmp[14] ),
    .S(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_1 _0968_ (.A(_0457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _0969_ (.A0(\SRAMController_ins.sram_data_out[15] ),
    .A1(\SRAMController_ins.sram_tmp[15] ),
    .S(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_1 _0970_ (.A(_0458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _0971_ (.A0(\SRAMController_ins.sram_data_out[16] ),
    .A1(\SRAMController_ins.sram_tmp[16] ),
    .S(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_1 _0972_ (.A(_0459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _0973_ (.A0(\SRAMController_ins.sram_data_out[17] ),
    .A1(\SRAMController_ins.sram_tmp[17] ),
    .S(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_1 _0974_ (.A(_0460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _0975_ (.A0(\SRAMController_ins.sram_data_out[18] ),
    .A1(\SRAMController_ins.sram_tmp[18] ),
    .S(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _0976_ (.A(_0461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _0977_ (.A0(\SRAMController_ins.sram_data_out[19] ),
    .A1(\SRAMController_ins.sram_tmp[19] ),
    .S(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_1 _0978_ (.A(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_4 _0979_ (.A(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _0980_ (.A0(\SRAMController_ins.sram_data_out[20] ),
    .A1(\SRAMController_ins.sram_tmp[20] ),
    .S(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0464_));
 sky130_fd_sc_hd__clkbuf_1 _0981_ (.A(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _0982_ (.A0(\SRAMController_ins.sram_data_out[21] ),
    .A1(\SRAMController_ins.sram_tmp[21] ),
    .S(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_1 _0983_ (.A(_0465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _0984_ (.A0(\SRAMController_ins.sram_data_out[22] ),
    .A1(\SRAMController_ins.sram_tmp[22] ),
    .S(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_1 _0985_ (.A(_0466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _0986_ (.A0(\SRAMController_ins.sram_data_out[23] ),
    .A1(\SRAMController_ins.sram_tmp[23] ),
    .S(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_1 _0987_ (.A(_0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _0988_ (.A0(\SRAMController_ins.sram_data_out[24] ),
    .A1(\SRAMController_ins.sram_tmp[24] ),
    .S(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_1 _0989_ (.A(_0468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _0990_ (.A0(\SRAMController_ins.sram_data_out[25] ),
    .A1(\SRAMController_ins.sram_tmp[25] ),
    .S(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_1 _0991_ (.A(_0469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _0992_ (.A0(\SRAMController_ins.sram_data_out[26] ),
    .A1(\SRAMController_ins.sram_tmp[26] ),
    .S(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0470_));
 sky130_fd_sc_hd__clkbuf_1 _0993_ (.A(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _0994_ (.A0(\SRAMController_ins.sram_data_out[27] ),
    .A1(\SRAMController_ins.sram_tmp[27] ),
    .S(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0471_));
 sky130_fd_sc_hd__clkbuf_1 _0995_ (.A(_0471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(\SRAMController_ins.sram_data_out[28] ),
    .A1(\SRAMController_ins.sram_tmp[28] ),
    .S(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_1 _0997_ (.A(_0472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _0998_ (.A0(\SRAMController_ins.sram_data_out[29] ),
    .A1(\SRAMController_ins.sram_tmp[29] ),
    .S(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_1 _0999_ (.A(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _1000_ (.A0(\SRAMController_ins.sram_data_out[30] ),
    .A1(\SRAMController_ins.sram_tmp[30] ),
    .S(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0474_));
 sky130_fd_sc_hd__clkbuf_1 _1001_ (.A(_0474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _1002_ (.A0(\SRAMController_ins.sram_data_out[31] ),
    .A1(\SRAMController_ins.sram_tmp[31] ),
    .S(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_1 _1003_ (.A(_0475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0106_));
 sky130_fd_sc_hd__and2_2 _1004_ (.A(\SRAMController_ins.rx_valid ),
    .B(_0236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0476_));
 sky130_fd_sc_hd__clkbuf_4 _1005_ (.A(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _1006_ (.A0(\SRAMController_ins.data_tmp[0] ),
    .A1(\SRAMController_ins.data_tmp[8] ),
    .S(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_1 _1007_ (.A(_0478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _1008_ (.A0(\SRAMController_ins.data_tmp[1] ),
    .A1(\SRAMController_ins.data_tmp[9] ),
    .S(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_1 _1009_ (.A(_0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _1010_ (.A0(\SRAMController_ins.data_tmp[2] ),
    .A1(\SRAMController_ins.data_tmp[10] ),
    .S(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0480_));
 sky130_fd_sc_hd__clkbuf_1 _1011_ (.A(_0480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _1012_ (.A0(\SRAMController_ins.data_tmp[3] ),
    .A1(\SRAMController_ins.data_tmp[11] ),
    .S(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0481_));
 sky130_fd_sc_hd__clkbuf_1 _1013_ (.A(_0481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _1014_ (.A0(\SRAMController_ins.data_tmp[4] ),
    .A1(\SRAMController_ins.data_tmp[12] ),
    .S(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0482_));
 sky130_fd_sc_hd__clkbuf_1 _1015_ (.A(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _1016_ (.A0(\SRAMController_ins.data_tmp[5] ),
    .A1(\SRAMController_ins.data_tmp[13] ),
    .S(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0483_));
 sky130_fd_sc_hd__clkbuf_1 _1017_ (.A(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _1018_ (.A0(\SRAMController_ins.data_tmp[6] ),
    .A1(\SRAMController_ins.data_tmp[14] ),
    .S(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0484_));
 sky130_fd_sc_hd__clkbuf_1 _1019_ (.A(_0484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _1020_ (.A0(\SRAMController_ins.data_tmp[7] ),
    .A1(\SRAMController_ins.data_tmp[15] ),
    .S(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_1 _1021_ (.A(_0485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _1022_ (.A0(\SRAMController_ins.data_tmp[8] ),
    .A1(\SRAMController_ins.data_tmp[16] ),
    .S(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0486_));
 sky130_fd_sc_hd__clkbuf_1 _1023_ (.A(_0486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _1024_ (.A0(\SRAMController_ins.data_tmp[9] ),
    .A1(\SRAMController_ins.data_tmp[17] ),
    .S(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_1 _1025_ (.A(_0487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_4 _1026_ (.A(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _1027_ (.A0(\SRAMController_ins.data_tmp[10] ),
    .A1(\SRAMController_ins.data_tmp[18] ),
    .S(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0489_));
 sky130_fd_sc_hd__clkbuf_1 _1028_ (.A(_0489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _1029_ (.A0(\SRAMController_ins.data_tmp[11] ),
    .A1(\SRAMController_ins.data_tmp[19] ),
    .S(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0490_));
 sky130_fd_sc_hd__clkbuf_1 _1030_ (.A(_0490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _1031_ (.A0(\SRAMController_ins.data_tmp[12] ),
    .A1(\SRAMController_ins.data_tmp[20] ),
    .S(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0491_));
 sky130_fd_sc_hd__clkbuf_1 _1032_ (.A(_0491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _1033_ (.A0(\SRAMController_ins.data_tmp[13] ),
    .A1(\SRAMController_ins.data_tmp[21] ),
    .S(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0492_));
 sky130_fd_sc_hd__clkbuf_1 _1034_ (.A(_0492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _1035_ (.A0(\SRAMController_ins.data_tmp[14] ),
    .A1(\SRAMController_ins.data_tmp[22] ),
    .S(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0493_));
 sky130_fd_sc_hd__clkbuf_1 _1036_ (.A(_0493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _1037_ (.A0(\SRAMController_ins.data_tmp[15] ),
    .A1(\SRAMController_ins.data_tmp[23] ),
    .S(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0494_));
 sky130_fd_sc_hd__clkbuf_1 _1038_ (.A(_0494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _1039_ (.A0(\SRAMController_ins.data_tmp[16] ),
    .A1(\SRAMController_ins.data_tmp[24] ),
    .S(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_1 _1040_ (.A(_0495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _1041_ (.A0(\SRAMController_ins.data_tmp[17] ),
    .A1(\SRAMController_ins.data_tmp[25] ),
    .S(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0496_));
 sky130_fd_sc_hd__clkbuf_1 _1042_ (.A(_0496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _1043_ (.A0(\SRAMController_ins.data_tmp[18] ),
    .A1(\SRAMController_ins.data_tmp[26] ),
    .S(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0497_));
 sky130_fd_sc_hd__clkbuf_1 _1044_ (.A(_0497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _1045_ (.A0(\SRAMController_ins.data_tmp[19] ),
    .A1(\SRAMController_ins.data_tmp[27] ),
    .S(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_1 _1046_ (.A(_0498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0126_));
 sky130_fd_sc_hd__clkbuf_4 _1047_ (.A(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _1048_ (.A0(\SRAMController_ins.data_tmp[20] ),
    .A1(\SRAMController_ins.data_tmp[28] ),
    .S(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0500_));
 sky130_fd_sc_hd__clkbuf_1 _1049_ (.A(_0500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _1050_ (.A0(\SRAMController_ins.data_tmp[21] ),
    .A1(\SRAMController_ins.data_tmp[29] ),
    .S(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_1 _1051_ (.A(_0501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _1052_ (.A0(\SRAMController_ins.data_tmp[22] ),
    .A1(\SRAMController_ins.data_tmp[30] ),
    .S(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0502_));
 sky130_fd_sc_hd__clkbuf_1 _1053_ (.A(_0502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _1054_ (.A0(\SRAMController_ins.data_tmp[23] ),
    .A1(\SRAMController_ins.data_tmp[31] ),
    .S(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0503_));
 sky130_fd_sc_hd__clkbuf_1 _1055_ (.A(_0503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _1056_ (.A0(\SRAMController_ins.data_tmp[24] ),
    .A1(\SRAMController_ins.rx_data_out[0] ),
    .S(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0504_));
 sky130_fd_sc_hd__clkbuf_1 _1057_ (.A(_0504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _1058_ (.A0(\SRAMController_ins.data_tmp[25] ),
    .A1(\SRAMController_ins.rx_data_out[1] ),
    .S(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0505_));
 sky130_fd_sc_hd__clkbuf_1 _1059_ (.A(_0505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _1060_ (.A0(\SRAMController_ins.data_tmp[26] ),
    .A1(\SRAMController_ins.rx_data_out[2] ),
    .S(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0506_));
 sky130_fd_sc_hd__clkbuf_1 _1061_ (.A(_0506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _1062_ (.A0(\SRAMController_ins.data_tmp[27] ),
    .A1(\SRAMController_ins.rx_data_out[3] ),
    .S(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0507_));
 sky130_fd_sc_hd__clkbuf_1 _1063_ (.A(_0507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _1064_ (.A0(\SRAMController_ins.data_tmp[28] ),
    .A1(\SRAMController_ins.rx_data_out[4] ),
    .S(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0508_));
 sky130_fd_sc_hd__clkbuf_1 _1065_ (.A(_0508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _1066_ (.A0(\SRAMController_ins.data_tmp[29] ),
    .A1(\SRAMController_ins.rx_data_out[5] ),
    .S(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0509_));
 sky130_fd_sc_hd__clkbuf_1 _1067_ (.A(_0509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _1068_ (.A0(\SRAMController_ins.data_tmp[30] ),
    .A1(\SRAMController_ins.rx_data_out[6] ),
    .S(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0510_));
 sky130_fd_sc_hd__clkbuf_1 _1069_ (.A(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _1070_ (.A0(\SRAMController_ins.data_tmp[31] ),
    .A1(\SRAMController_ins.rx_data_out[7] ),
    .S(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0511_));
 sky130_fd_sc_hd__clkbuf_1 _1071_ (.A(_0511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(_0138_));
 sky130_fd_sc_hd__dfxtp_1 _1072_ (.CLK(clknet_4_6_0_clk),
    .D(_0008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.out_latched ));
 sky130_fd_sc_hd__dfxtp_1 _1073_ (.CLK(clknet_4_5_0_clk),
    .D(_0009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1074_ (.CLK(clknet_4_5_0_clk),
    .D(_0010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1075_ (.CLK(clknet_4_5_0_clk),
    .D(_0011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1076_ (.CLK(clknet_4_5_0_clk),
    .D(_0012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1077_ (.CLK(clknet_4_5_0_clk),
    .D(_0013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1078_ (.CLK(clknet_4_5_0_clk),
    .D(_0014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1079_ (.CLK(clknet_4_5_0_clk),
    .D(_0015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.CLK(clknet_4_6_0_clk),
    .D(_0016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.data[7] ));
 sky130_fd_sc_hd__dfxtp_2 _1081_ (.CLK(clknet_4_7_0_clk),
    .D(_0017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.sampleCount[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1082_ (.CLK(clknet_4_7_0_clk),
    .D(_0018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.sampleCount[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1083_ (.CLK(clknet_4_7_0_clk),
    .D(_0019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.sampleCount[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1084_ (.CLK(clknet_4_6_0_clk),
    .D(_0020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.sampleCount[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1085_ (.CLK(clknet_4_6_0_clk),
    .D(_0021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.inputReg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.CLK(clknet_4_7_0_clk),
    .D(_0022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.inputReg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1087_ (.CLK(clknet_4_7_0_clk),
    .D(_0023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.inputReg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1088_ (.CLK(clknet_4_5_0_clk),
    .D(_0024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.bitIndex[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1089_ (.CLK(clknet_4_5_0_clk),
    .D(_0025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.bitIndex[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1090_ (.CLK(clknet_4_5_0_clk),
    .D(_0026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.bitIndex[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1091_ (.CLK(clknet_4_4_0_clk),
    .D(_0027_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.addr_tmp[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1092_ (.CLK(clknet_4_4_0_clk),
    .D(_0028_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.addr_tmp[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1093_ (.CLK(clknet_4_4_0_clk),
    .D(_0029_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.addr_tmp[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1094_ (.CLK(clknet_4_4_0_clk),
    .D(_0030_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.addr_tmp[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1095_ (.CLK(clknet_4_5_0_clk),
    .D(_0031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.overrun ));
 sky130_fd_sc_hd__dfxtp_1 _1096_ (.CLK(clknet_4_5_0_clk),
    .D(_0032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.error ));
 sky130_fd_sc_hd__dfxtp_2 _1097_ (.CLK(clknet_4_13_0_clk),
    .D(_0033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_valid ));
 sky130_fd_sc_hd__dfxtp_1 _1098_ (.CLK(clknet_4_4_0_clk),
    .D(_0034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1099_ (.CLK(clknet_4_4_0_clk),
    .D(_0035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1100_ (.CLK(clknet_4_5_0_clk),
    .D(_0036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1101_ (.CLK(clknet_4_4_0_clk),
    .D(_0037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1102_ (.CLK(clknet_4_4_0_clk),
    .D(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[4] ));
 sky130_fd_sc_hd__dfxtp_2 _1103_ (.CLK(clknet_4_5_0_clk),
    .D(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1104_ (.CLK(clknet_4_4_0_clk),
    .D(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1105_ (.CLK(clknet_4_4_0_clk),
    .D(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.rx_data_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1106_ (.CLK(clknet_4_9_0_clk),
    .D(_0042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1107_ (.CLK(clknet_4_14_0_clk),
    .D(_0043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1108_ (.CLK(clknet_4_9_0_clk),
    .D(_0044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1109_ (.CLK(clknet_4_8_0_clk),
    .D(_0045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1110_ (.CLK(clknet_4_8_0_clk),
    .D(_0046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1111_ (.CLK(clknet_4_8_0_clk),
    .D(_0047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1112_ (.CLK(clknet_4_9_0_clk),
    .D(_0048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1113_ (.CLK(clknet_4_9_0_clk),
    .D(_0049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1114_ (.CLK(clknet_4_9_0_clk),
    .D(_0050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1115_ (.CLK(clknet_4_14_0_clk),
    .D(_0051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1116_ (.CLK(clknet_4_14_0_clk),
    .D(_0052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1117_ (.CLK(clknet_4_14_0_clk),
    .D(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.txCounter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1118_ (.CLK(clknet_4_12_0_clk),
    .D(_0054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1119_ (.CLK(clknet_4_12_0_clk),
    .D(_0055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1120_ (.CLK(clknet_4_12_0_clk),
    .D(_0056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1121_ (.CLK(clknet_4_12_0_clk),
    .D(_0057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1122_ (.CLK(clknet_4_15_0_clk),
    .D(_0058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1123_ (.CLK(clknet_4_15_0_clk),
    .D(_0059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1124_ (.CLK(clknet_4_12_0_clk),
    .D(_0060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1125_ (.CLK(clknet_4_12_0_clk),
    .D(_0061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.data[7] ));
 sky130_fd_sc_hd__dfxtp_2 _1126_ (.CLK(clknet_4_14_0_clk),
    .D(_0062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.bitIndex[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1127_ (.CLK(clknet_4_9_0_clk),
    .D(_0063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.bitIndex[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1128_ (.CLK(clknet_4_15_0_clk),
    .D(_0064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.bitIndex[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1129_ (.CLK(clknet_4_15_0_clk),
    .D(_0065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.out ));
 sky130_fd_sc_hd__dfxtp_1 _1130_ (.CLK(clknet_4_15_0_clk),
    .D(_0066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.tx_ready ));
 sky130_fd_sc_hd__dfxtp_1 _1131_ (.CLK(clknet_4_15_0_clk),
    .D(_0004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1132_ (.CLK(clknet_4_15_0_clk),
    .D(_0005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1133_ (.CLK(clknet_4_14_0_clk),
    .D(_0006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1134_ (.CLK(clknet_4_15_0_clk),
    .D(_0007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTTransmitter_ins.state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1135_ (.CLK(clknet_4_7_0_clk),
    .D(_0067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1136_ (.CLK(clknet_4_13_0_clk),
    .D(_0068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1137_ (.CLK(clknet_4_13_0_clk),
    .D(_0069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1138_ (.CLK(clknet_4_13_0_clk),
    .D(_0070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1139_ (.CLK(clknet_4_7_0_clk),
    .D(_0071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1140_ (.CLK(clknet_4_7_0_clk),
    .D(_0072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[5] ));
 sky130_fd_sc_hd__dfxtp_4 _1141_ (.CLK(clknet_4_13_0_clk),
    .D(_0073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[6] ));
 sky130_fd_sc_hd__dfxtp_4 _1142_ (.CLK(clknet_4_13_0_clk),
    .D(_0074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.rxCounter[7] ));
 sky130_fd_sc_hd__dfxtp_2 _1143_ (.CLK(clknet_4_7_0_clk),
    .D(_0000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1144_ (.CLK(clknet_4_6_0_clk),
    .D(_0001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1145_ (.CLK(clknet_4_6_0_clk),
    .D(_0002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1146_ (.CLK(clknet_4_6_0_clk),
    .D(_0003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\UARTReceiver_ins.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1147_ (.CLK(clknet_4_3_0_clk),
    .D(_0075_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1148_ (.CLK(clknet_4_13_0_clk),
    .D(_0076_),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1149_ (.CLK(clknet_4_2_0_clk),
    .D(_0077_),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1150_ (.CLK(clknet_4_0_0_clk),
    .D(_0078_),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1151_ (.CLK(clknet_4_2_0_clk),
    .D(_0079_),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[4] ));
 sky130_fd_sc_hd__dfrtp_4 _1152_ (.CLK(clknet_4_2_0_clk),
    .D(_0080_),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1153_ (.CLK(clknet_4_2_0_clk),
    .D(_0081_),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[6] ));
 sky130_fd_sc_hd__dfrtp_2 _1154_ (.CLK(clknet_4_2_0_clk),
    .D(_0082_),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1155_ (.CLK(clknet_4_0_0_clk),
    .D(_0083_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1156_ (.CLK(clknet_4_12_0_clk),
    .D(_0084_),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1157_ (.CLK(clknet_4_3_0_clk),
    .D(_0085_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1158_ (.CLK(clknet_4_2_0_clk),
    .D(_0086_),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1159_ (.CLK(clknet_4_8_0_clk),
    .D(_0087_),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1160_ (.CLK(clknet_4_11_0_clk),
    .D(_0088_),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1161_ (.CLK(clknet_4_12_0_clk),
    .D(_0089_),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1162_ (.CLK(clknet_4_10_0_clk),
    .D(_0090_),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1163_ (.CLK(clknet_4_3_0_clk),
    .D(_0091_),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1164_ (.CLK(clknet_4_13_0_clk),
    .D(_0092_),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1165_ (.CLK(clknet_4_3_0_clk),
    .D(_0093_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1166_ (.CLK(clknet_4_2_0_clk),
    .D(_0094_),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[19] ));
 sky130_fd_sc_hd__dfrtp_2 _1167_ (.CLK(clknet_4_11_0_clk),
    .D(_0095_),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[20] ));
 sky130_fd_sc_hd__dfrtp_2 _1168_ (.CLK(clknet_4_11_0_clk),
    .D(_0096_),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[21] ));
 sky130_fd_sc_hd__dfrtp_4 _1169_ (.CLK(clknet_4_11_0_clk),
    .D(_0097_),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[22] ));
 sky130_fd_sc_hd__dfrtp_2 _1170_ (.CLK(clknet_4_11_0_clk),
    .D(_0098_),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[23] ));
 sky130_fd_sc_hd__dfrtp_4 _1171_ (.CLK(clknet_4_10_0_clk),
    .D(_0099_),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[24] ));
 sky130_fd_sc_hd__dfrtp_4 _1172_ (.CLK(clknet_4_10_0_clk),
    .D(_0100_),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[25] ));
 sky130_fd_sc_hd__dfrtp_4 _1173_ (.CLK(clknet_4_10_0_clk),
    .D(_0101_),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[26] ));
 sky130_fd_sc_hd__dfrtp_4 _1174_ (.CLK(clknet_4_10_0_clk),
    .D(_0102_),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[27] ));
 sky130_fd_sc_hd__dfrtp_1 _1175_ (.CLK(clknet_4_10_0_clk),
    .D(_0103_),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[28] ));
 sky130_fd_sc_hd__dfrtp_1 _1176_ (.CLK(clknet_4_11_0_clk),
    .D(_0104_),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[29] ));
 sky130_fd_sc_hd__dfrtp_4 _1177_ (.CLK(clknet_4_11_0_clk),
    .D(_0105_),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1178_ (.CLK(clknet_4_11_0_clk),
    .D(_0106_),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.sram_tmp[31] ));
 sky130_fd_sc_hd__dfrtp_4 _1179_ (.CLK(clknet_4_13_0_clk),
    .D(\SRAMController_ins.nxt_state[0] ),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.cur_state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1180_ (.CLK(clknet_4_13_0_clk),
    .D(\SRAMController_ins.nxt_state[1] ),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.cur_state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1181_ (.CLK(clknet_4_13_0_clk),
    .D(\SRAMController_ins.nxt_state[2] ),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.cur_state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1182_ (.CLK(clknet_4_13_0_clk),
    .D(\SRAMController_ins.nxt_state[3] ),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.cur_state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1183_ (.CLK(clknet_4_3_0_clk),
    .D(_0107_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1184_ (.CLK(clknet_4_3_0_clk),
    .D(_0108_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1185_ (.CLK(clknet_4_3_0_clk),
    .D(_0109_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1186_ (.CLK(clknet_4_3_0_clk),
    .D(_0110_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1187_ (.CLK(clknet_4_0_0_clk),
    .D(_0111_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1188_ (.CLK(clknet_4_3_0_clk),
    .D(_0112_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1189_ (.CLK(clknet_4_0_0_clk),
    .D(_0113_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1190_ (.CLK(clknet_4_3_0_clk),
    .D(_0114_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1191_ (.CLK(clknet_4_3_0_clk),
    .D(_0115_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1192_ (.CLK(clknet_4_0_0_clk),
    .D(_0116_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1193_ (.CLK(clknet_4_3_0_clk),
    .D(_0117_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1194_ (.CLK(clknet_4_3_0_clk),
    .D(_0118_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1195_ (.CLK(clknet_4_0_0_clk),
    .D(_0119_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1196_ (.CLK(clknet_4_3_0_clk),
    .D(_0120_),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1197_ (.CLK(clknet_4_0_0_clk),
    .D(_0121_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1198_ (.CLK(clknet_4_3_0_clk),
    .D(_0122_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1199_ (.CLK(clknet_4_2_0_clk),
    .D(_0123_),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1200_ (.CLK(clknet_4_2_0_clk),
    .D(_0124_),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1201_ (.CLK(clknet_4_0_0_clk),
    .D(_0125_),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1202_ (.CLK(clknet_4_0_0_clk),
    .D(_0126_),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[19] ));
 sky130_fd_sc_hd__dfrtp_1 _1203_ (.CLK(clknet_4_0_0_clk),
    .D(_0127_),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1204_ (.CLK(clknet_4_0_0_clk),
    .D(_0128_),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1205_ (.CLK(clknet_4_0_0_clk),
    .D(_0129_),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1206_ (.CLK(clknet_4_1_0_clk),
    .D(_0130_),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[23] ));
 sky130_fd_sc_hd__dfrtp_1 _1207_ (.CLK(clknet_4_1_0_clk),
    .D(_0131_),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[24] ));
 sky130_fd_sc_hd__dfrtp_1 _1208_ (.CLK(clknet_4_1_0_clk),
    .D(_0132_),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[25] ));
 sky130_fd_sc_hd__dfrtp_1 _1209_ (.CLK(clknet_4_1_0_clk),
    .D(_0133_),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[26] ));
 sky130_fd_sc_hd__dfrtp_1 _1210_ (.CLK(clknet_4_1_0_clk),
    .D(_0134_),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[27] ));
 sky130_fd_sc_hd__dfrtp_1 _1211_ (.CLK(clknet_4_1_0_clk),
    .D(_0135_),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[28] ));
 sky130_fd_sc_hd__dfrtp_1 _1212_ (.CLK(clknet_4_1_0_clk),
    .D(_0136_),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[29] ));
 sky130_fd_sc_hd__dfrtp_1 _1213_ (.CLK(clknet_4_1_0_clk),
    .D(_0137_),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1214_ (.CLK(clknet_4_1_0_clk),
    .D(_0138_),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .Q(\SRAMController_ins.data_tmp[31] ));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .HI(net56));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__conb_1 sram_ins_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net31));
 sky130_fd_sc_hd__conb_1 sram_ins_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net32));
 sky130_fd_sc_hd__conb_1 sram_ins_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net33));
 sky130_fd_sc_hd__conb_1 sram_ins_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net34));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net35));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net36));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net37));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net38));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net39));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net40));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net41));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net42));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net43));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net44));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net45));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net46));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net47));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net48));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net49));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net50));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net51));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net52));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net53));
 sky130_fd_sc_hd__conb_1 tt_um_kmakise_sram_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net54));
 sky130_fd_sc_hd__conb_1 sram_ins_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .HI(net55));
 sky130_fd_sc_hd__buf_4 _1242_ (.A(\UARTTransmitter_ins.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(uio_out[4]));
 sky130_fd_sc_hd__clkbuf_4 _1243_ (.A(\UARTReceiver_ins.overrun ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__clkbuf_4 _1244_ (.A(\UARTReceiver_ins.error ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(uo_out[7]));
 myconfig_sky_dual sram_ins (.csb0(\SRAMController_ins.csb_n ),
    .csb1(net55),
    .web0(\SRAMController_ins.we_n ),
    .clk0(clknet_4_2_0_clk),
    .clk1(net34),
    .vccd1(VDPWR),
    .vssd1(VGND),
    .addr0({\SRAMController_ins.addr[3] ,
    \SRAMController_ins.addr[2] ,
    \SRAMController_ins.addr[1] ,
    \SRAMController_ins.addr[0] }),
    .addr1({net33,
    net32,
    net31,
    net30}),
    .din0({\SRAMController_ins.sram_data_in[31] ,
    \SRAMController_ins.sram_data_in[30] ,
    \SRAMController_ins.sram_data_in[29] ,
    \SRAMController_ins.sram_data_in[28] ,
    \SRAMController_ins.sram_data_in[27] ,
    \SRAMController_ins.sram_data_in[26] ,
    \SRAMController_ins.sram_data_in[25] ,
    \SRAMController_ins.sram_data_in[24] ,
    \SRAMController_ins.sram_data_in[23] ,
    \SRAMController_ins.sram_data_in[22] ,
    \SRAMController_ins.sram_data_in[21] ,
    \SRAMController_ins.sram_data_in[20] ,
    \SRAMController_ins.sram_data_in[19] ,
    \SRAMController_ins.sram_data_in[18] ,
    \SRAMController_ins.sram_data_in[17] ,
    \SRAMController_ins.sram_data_in[16] ,
    \SRAMController_ins.sram_data_in[15] ,
    \SRAMController_ins.sram_data_in[14] ,
    \SRAMController_ins.sram_data_in[13] ,
    \SRAMController_ins.sram_data_in[12] ,
    \SRAMController_ins.sram_data_in[11] ,
    \SRAMController_ins.sram_data_in[10] ,
    \SRAMController_ins.sram_data_in[9] ,
    \SRAMController_ins.sram_data_in[8] ,
    \SRAMController_ins.sram_data_in[7] ,
    \SRAMController_ins.sram_data_in[6] ,
    \SRAMController_ins.sram_data_in[5] ,
    \SRAMController_ins.sram_data_in[4] ,
    \SRAMController_ins.sram_data_in[3] ,
    \SRAMController_ins.sram_data_in[2] ,
    \SRAMController_ins.sram_data_in[1] ,
    \SRAMController_ins.sram_data_in[0] }),
    .dout0({\SRAMController_ins.sram_data_out[31] ,
    \SRAMController_ins.sram_data_out[30] ,
    \SRAMController_ins.sram_data_out[29] ,
    \SRAMController_ins.sram_data_out[28] ,
    \SRAMController_ins.sram_data_out[27] ,
    \SRAMController_ins.sram_data_out[26] ,
    \SRAMController_ins.sram_data_out[25] ,
    \SRAMController_ins.sram_data_out[24] ,
    \SRAMController_ins.sram_data_out[23] ,
    \SRAMController_ins.sram_data_out[22] ,
    \SRAMController_ins.sram_data_out[21] ,
    \SRAMController_ins.sram_data_out[20] ,
    \SRAMController_ins.sram_data_out[19] ,
    \SRAMController_ins.sram_data_out[18] ,
    \SRAMController_ins.sram_data_out[17] ,
    \SRAMController_ins.sram_data_out[16] ,
    \SRAMController_ins.sram_data_out[15] ,
    \SRAMController_ins.sram_data_out[14] ,
    \SRAMController_ins.sram_data_out[13] ,
    \SRAMController_ins.sram_data_out[12] ,
    \SRAMController_ins.sram_data_out[11] ,
    \SRAMController_ins.sram_data_out[10] ,
    \SRAMController_ins.sram_data_out[9] ,
    \SRAMController_ins.sram_data_out[8] ,
    \SRAMController_ins.sram_data_out[7] ,
    \SRAMController_ins.sram_data_out[6] ,
    \SRAMController_ins.sram_data_out[5] ,
    \SRAMController_ins.sram_data_out[4] ,
    \SRAMController_ins.sram_data_out[3] ,
    \SRAMController_ins.sram_data_out[2] ,
    \SRAMController_ins.sram_data_out[1] ,
    \SRAMController_ins.sram_data_out[0] }),
    .dout1({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16,
    _NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32}));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_2_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_2_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_2_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_2_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_2_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_2_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_2_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_2_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_2_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Right_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Right_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Right_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Right_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Right_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Right_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Right_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Right_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Right_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Right_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Right_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Right_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Right_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Right_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Right_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Right_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Right_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Right_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Right_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Right_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Right_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Right_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Right_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Right_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Right_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Right_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Right_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Right_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Right_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Right_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Right_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Right_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Right_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Right_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Right_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Right_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Right_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Right_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Right_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Right_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Right_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Right_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_1_Left_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_1_Left_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_1_Left_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_1_Left_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_1_Left_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_1_Left_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_1_Left_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_1_Left_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Left_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Left_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Left_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Left_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Left_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Left_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Left_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Left_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Left_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Left_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Left_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Left_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Left_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Left_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Left_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Left_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Left_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Left_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Left_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Left_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Left_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Left_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Left_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Left_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Left_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Left_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Left_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Left_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Left_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Left_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Left_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Left_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Left_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Left_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Left_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Left_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Left_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Left_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Left_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Left_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Left_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Left_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Left_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Left_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Left_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Left_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Left_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Left_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Left_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Left_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Left_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Left_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Left_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Left_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Left_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Left_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Left_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Left_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Left_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Left_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_1_Left_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_2_Left_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_2_Left_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_2_Left_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_2_Left_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_2_Left_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_2_Left_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_2_Left_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_2_Left_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_2_Left_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Left_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Left_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Left_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Left_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Left_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Left_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Left_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Left_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Left_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Left_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Left_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Left_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Left_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Left_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Left_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Left_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Left_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Left_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Left_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Left_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Left_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Left_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Left_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Left_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Left_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Left_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Left_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Left_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Left_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Left_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Left_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Left_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Left_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Left_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Left_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Left_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Left_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Left_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Left_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Left_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Left_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Left_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Left_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Left_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Left_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Left_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Left_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Left_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Left_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Left_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Left_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Left_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Left_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Left_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Left_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Left_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Left_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Left_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Left_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Left_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_1_Right_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_1_Right_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_1_Right_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_1_Right_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_1_Right_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_1_Right_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_1_Right_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_1_Right_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Right_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Right_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Right_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Right_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Right_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Right_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Right_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Right_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Right_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Right_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Right_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Right_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Right_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Right_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Right_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Right_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Right_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Right_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Right_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Right_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Right_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Right_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Right_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Right_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Right_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Right_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Right_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Right_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Right_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Right_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Right_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Right_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Right_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Right_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Right_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Right_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Right_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Right_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Right_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Right_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Right_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Right_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Right_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Right_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Right_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Right_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Right_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Right_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Right_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Right_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Right_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Right_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Right_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Right_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Right_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Right_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Right_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Right_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Right_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Right_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_1_Right_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_300 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_301 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_302 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_303 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_304 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_305 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_306 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_307 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_308 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_309 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_310 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_311 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_312 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_313 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_314 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_315 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_316 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_317 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_318 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_319 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_320 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_321 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_322 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_323 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_324 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_325 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_326 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_327 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_328 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_329 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_330 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_331 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_332 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_333 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_334 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_335 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_336 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_337 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1_338 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1_339 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1_340 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1_341 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1_342 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1_343 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1_344 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1_345 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1_346 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1_347 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1_348 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1_349 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1_350 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1_351 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1_352 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1_353 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1_354 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1_355 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1_356 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1_357 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1_358 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1_359 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1_360 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1_361 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_1_362 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_1_363 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_1_364 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_1_365 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_1_366 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_1_367 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_1_368 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_1_369 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_1_370 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_1_371 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_1_372 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_1_373 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1_374 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1_375 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1_376 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1_377 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1_378 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1_379 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1_380 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1_381 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1_382 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1_383 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1_384 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1_385 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1_386 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1_387 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1_388 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1_389 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1_390 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1_391 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1_392 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1_393 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1_394 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1_395 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1_396 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1_397 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1_398 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1_399 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1_400 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1_401 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1_402 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1_403 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1_404 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1_405 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1_406 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1_407 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1_408 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1_409 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1_410 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1_411 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1_412 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1_413 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1_414 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1_415 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1_416 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1_417 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1_418 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1_419 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1_420 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1_421 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1_422 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1_423 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1_424 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1_425 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1_426 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1_427 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1_428 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1_429 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1_430 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1_431 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1_432 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1_433 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1_434 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1_435 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1_436 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1_437 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1_438 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1_439 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1_440 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1_441 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1_442 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1_443 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1_444 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1_445 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1_446 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1_447 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1_448 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1_449 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1_450 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1_451 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1_452 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1_453 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1_454 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1_455 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1_456 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1_457 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1_458 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1_459 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1_460 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1_461 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1_462 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1_463 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1_464 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1_465 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1_466 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1_467 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1_468 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1_469 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1_470 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1_471 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1_472 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1_473 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1_474 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1_475 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1_476 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1_477 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1_478 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1_479 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1_480 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1_481 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1_482 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1_483 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1_484 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1_485 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1_486 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1_487 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1_488 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1_489 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1_490 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1_491 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1_492 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1_493 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1_494 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1_495 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1_496 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1_497 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1_498 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1_499 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1_500 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1_501 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1_502 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1_503 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1_504 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1_505 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1_506 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1_507 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1_508 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1_509 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1_510 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1_511 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1_512 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1_513 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1_514 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1_515 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1_516 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1_517 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1_518 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1_519 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1_520 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1_521 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1_522 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1_523 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1_524 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1_525 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1_526 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1_527 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1_528 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1_529 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1_530 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1_531 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1_532 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1_533 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1_534 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1_535 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1_536 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1_537 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1_538 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1_539 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1_540 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1_541 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_542 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_543 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_544 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_545 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_546 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_547 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_548 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_549 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_550 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_551 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_552 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_553 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_554 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_555 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_556 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_557 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_558 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_559 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_560 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_561 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_562 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_563 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_564 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_565 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_566 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_567 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_568 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_569 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_570 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_571 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_572 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_573 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_574 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_575 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_576 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_577 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_578 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_579 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_580 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_581 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_582 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_583 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_584 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_585 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_586 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_587 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_588 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_589 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_590 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_591 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_592 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_593 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_594 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_595 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_596 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_597 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_598 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_599 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_600 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_601 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_602 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_603 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_604 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_605 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_606 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_607 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_608 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_609 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_610 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_611 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_612 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_613 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_614 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_615 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_616 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_617 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_618 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_619 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_620 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_621 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_622 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_623 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_624 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_625 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_626 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_627 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_628 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_629 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_630 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_631 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_632 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_633 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_634 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_635 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_636 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_637 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_638 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_639 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_640 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_641 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_642 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_643 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_644 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_645 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_646 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_647 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_648 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_649 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_650 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_651 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_652 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_653 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_654 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_655 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_656 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_657 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_658 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_659 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_660 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_661 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_662 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_663 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_664 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_665 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_666 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_667 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_668 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_669 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_670 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_671 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_672 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_673 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_674 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_675 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_676 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_677 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_678 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_679 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_680 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_681 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_682 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_683 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_684 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_685 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_686 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_687 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_688 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_689 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_690 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_691 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_692 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_693 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_694 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_695 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_696 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_697 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_698 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_699 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_700 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_701 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_702 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_703 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_704 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_705 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_706 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_707 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_708 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_709 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_710 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_711 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_712 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_713 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_714 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_715 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_716 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_717 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_718 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_719 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_720 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_721 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_722 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_723 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_724 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_725 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_726 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_727 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_728 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_729 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_730 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_731 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_732 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_733 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_734 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_735 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_736 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_737 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_738 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_739 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_740 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_741 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_742 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_743 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_744 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_745 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_746 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_747 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_748 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_749 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_750 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_751 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_752 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_753 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_754 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_755 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_756 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_757 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_758 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_759 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_760 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_761 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_762 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_763 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_764 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_765 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_766 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_767 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_768 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_769 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_770 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_771 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_772 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_773 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_774 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_775 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_776 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_777 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_778 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_779 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_780 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_781 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_782 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_783 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_784 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_785 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_786 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_787 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_788 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1_789 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1_790 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1_791 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_2_792 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_2_793 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_2_794 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_2_795 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_2_796 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_2_797 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_2_798 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_2_799 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_2_800 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_801 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_2_802 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_803 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_2_804 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_805 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_2_806 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_807 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_2_808 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_809 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_2_810 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_811 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_2_812 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_813 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_2_814 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_815 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_2_816 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_817 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_2_818 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_819 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_2_820 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_821 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2_822 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_823 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2_824 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_825 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_2_826 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_827 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_2_828 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_829 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_2_830 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_831 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_2_832 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_833 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_2_834 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_835 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_2_836 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_837 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_2_838 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_839 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_2_840 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_841 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_2_842 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_843 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_2_844 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_845 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_2_846 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_847 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2_848 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_849 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2_850 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_851 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2_852 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_853 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2_854 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_855 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2_856 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_857 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2_858 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_859 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2_860 (.VGND(VGND),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 max_cap3 (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap4 (.A(_0176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 wire5 (.A(_0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 max_cap6 (.A(_0167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 max_cap7 (.A(_0166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net7));
 sky130_fd_sc_hd__buf_2 fanout8 (.A(\UARTReceiver_ins.state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 fanout9 (.A(\UARTReceiver_ins.state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net9));
 sky130_fd_sc_hd__buf_2 fanout10 (.A(\UARTReceiver_ins.state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net10));
 sky130_fd_sc_hd__buf_2 fanout11 (.A(\SRAMController_ins.tx_ready ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 fanout12 (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 fanout15 (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net15));
 sky130_fd_sc_hd__buf_2 fanout16 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout20 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 fanout22 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout23 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net23));
 sky130_fd_sc_hd__buf_2 fanout24 (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net24));
 sky130_fd_sc_hd__buf_1 fanout25 (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net25));
 sky130_fd_sc_hd__buf_2 fanout26 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net28));
 sky130_fd_sc_hd__buf_4 fanout29 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net29));
 sky130_fd_sc_hd__conb_1 sram_ins_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .LO(net30));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload0 (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__clkinv_4 clkload1 (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__clkinv_4 clkload2 (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_4 clkload3 (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload4 (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_6 clkload5 (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__clkinv_4 clkload6 (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__clkinv_8 clkload7 (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_8 clkload8 (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_8 clkload9 (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_6 clkload10 (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_6 clkload11 (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__clkinv_2 clkload12 (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_8 clkload13 (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__inv_6 clkload14 (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\UARTTransmitter_ins.txCounter[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\UARTTransmitter_ins.state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\UARTReceiver_ins.rxCounter[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\UARTReceiver_ins.data[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\UARTReceiver_ins.data[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\UARTTransmitter_ins.data[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\UARTTransmitter_ins.data[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\UARTTransmitter_ins.data[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\UARTTransmitter_ins.data[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\UARTReceiver_ins.data[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\UARTReceiver_ins.data[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\UARTTransmitter_ins.data[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\UARTReceiver_ins.inputReg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\UARTReceiver_ins.error ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\UARTReceiver_ins.data[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\UARTReceiver_ins.data[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\UARTReceiver_ins.data[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\UARTReceiver_ins.data[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\UARTReceiver_ins.inputReg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\UARTReceiver_ins.inputReg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\UARTReceiver_ins.state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\UARTReceiver_ins.rxCounter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\SRAMController_ins.rx_valid ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\UARTReceiver_ins.data[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR),
    .X(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1098__Q (.DIODE(\SRAMController_ins.rx_data_out[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1056__A1 (.DIODE(\SRAMController_ins.rx_data_out[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__A1 (.DIODE(\SRAMController_ins.rx_data_out[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__A1 (.DIODE(\SRAMController_ins.rx_data_out[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__B2 (.DIODE(\SRAMController_ins.rx_data_out[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1099__Q (.DIODE(\SRAMController_ins.rx_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1058__A1 (.DIODE(\SRAMController_ins.rx_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0795__A1 (.DIODE(\SRAMController_ins.rx_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__A1 (.DIODE(\SRAMController_ins.rx_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__B2 (.DIODE(\SRAMController_ins.rx_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1100__Q (.DIODE(\SRAMController_ins.rx_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1060__A1 (.DIODE(\SRAMController_ins.rx_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0796__A1 (.DIODE(\SRAMController_ins.rx_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__A1 (.DIODE(\SRAMController_ins.rx_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__B2 (.DIODE(\SRAMController_ins.rx_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1101__Q (.DIODE(\SRAMController_ins.rx_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1062__A1 (.DIODE(\SRAMController_ins.rx_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__A1 (.DIODE(\SRAMController_ins.rx_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__A1 (.DIODE(\SRAMController_ins.rx_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__B2 (.DIODE(\SRAMController_ins.rx_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__Q (.DIODE(\SRAMController_ins.rx_data_out[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1064__A1 (.DIODE(\SRAMController_ins.rx_data_out[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0798__A1 (.DIODE(\SRAMController_ins.rx_data_out[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1103__Q (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1066__A1 (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0799__A1 (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0666__A_N (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0651__A (.DIODE(\SRAMController_ins.rx_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[0]  (.DIODE(\SRAMController_ins.sram_data_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0585__X (.DIODE(\SRAMController_ins.sram_data_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[10]  (.DIODE(\SRAMController_ins.sram_data_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0606__X (.DIODE(\SRAMController_ins.sram_data_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[11]  (.DIODE(\SRAMController_ins.sram_data_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0608__X (.DIODE(\SRAMController_ins.sram_data_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[12]  (.DIODE(\SRAMController_ins.sram_data_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0610__X (.DIODE(\SRAMController_ins.sram_data_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[13]  (.DIODE(\SRAMController_ins.sram_data_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0612__X (.DIODE(\SRAMController_ins.sram_data_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[14]  (.DIODE(\SRAMController_ins.sram_data_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0614__X (.DIODE(\SRAMController_ins.sram_data_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[15]  (.DIODE(\SRAMController_ins.sram_data_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0617__X (.DIODE(\SRAMController_ins.sram_data_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[16]  (.DIODE(\SRAMController_ins.sram_data_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0619__X (.DIODE(\SRAMController_ins.sram_data_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[17]  (.DIODE(\SRAMController_ins.sram_data_in[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0621__X (.DIODE(\SRAMController_ins.sram_data_in[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[18]  (.DIODE(\SRAMController_ins.sram_data_in[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0623__X (.DIODE(\SRAMController_ins.sram_data_in[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[19]  (.DIODE(\SRAMController_ins.sram_data_in[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0625__X (.DIODE(\SRAMController_ins.sram_data_in[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[1]  (.DIODE(\SRAMController_ins.sram_data_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0587__X (.DIODE(\SRAMController_ins.sram_data_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[20]  (.DIODE(\SRAMController_ins.sram_data_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0627__X (.DIODE(\SRAMController_ins.sram_data_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[21]  (.DIODE(\SRAMController_ins.sram_data_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0629__X (.DIODE(\SRAMController_ins.sram_data_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[22]  (.DIODE(\SRAMController_ins.sram_data_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0631__X (.DIODE(\SRAMController_ins.sram_data_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[23]  (.DIODE(\SRAMController_ins.sram_data_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0633__X (.DIODE(\SRAMController_ins.sram_data_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[24]  (.DIODE(\SRAMController_ins.sram_data_in[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0635__X (.DIODE(\SRAMController_ins.sram_data_in[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[25]  (.DIODE(\SRAMController_ins.sram_data_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__X (.DIODE(\SRAMController_ins.sram_data_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[26]  (.DIODE(\SRAMController_ins.sram_data_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0639__X (.DIODE(\SRAMController_ins.sram_data_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[27]  (.DIODE(\SRAMController_ins.sram_data_in[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0641__X (.DIODE(\SRAMController_ins.sram_data_in[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[28]  (.DIODE(\SRAMController_ins.sram_data_in[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0643__X (.DIODE(\SRAMController_ins.sram_data_in[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[29]  (.DIODE(\SRAMController_ins.sram_data_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0645__X (.DIODE(\SRAMController_ins.sram_data_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[2]  (.DIODE(\SRAMController_ins.sram_data_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0589__X (.DIODE(\SRAMController_ins.sram_data_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[30]  (.DIODE(\SRAMController_ins.sram_data_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0647__X (.DIODE(\SRAMController_ins.sram_data_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[31]  (.DIODE(\SRAMController_ins.sram_data_in[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0649__X (.DIODE(\SRAMController_ins.sram_data_in[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[3]  (.DIODE(\SRAMController_ins.sram_data_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0591__X (.DIODE(\SRAMController_ins.sram_data_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[4]  (.DIODE(\SRAMController_ins.sram_data_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0593__X (.DIODE(\SRAMController_ins.sram_data_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[5]  (.DIODE(\SRAMController_ins.sram_data_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0596__X (.DIODE(\SRAMController_ins.sram_data_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[6]  (.DIODE(\SRAMController_ins.sram_data_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0598__X (.DIODE(\SRAMController_ins.sram_data_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[7]  (.DIODE(\SRAMController_ins.sram_data_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0600__X (.DIODE(\SRAMController_ins.sram_data_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[8]  (.DIODE(\SRAMController_ins.sram_data_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0602__X (.DIODE(\SRAMController_ins.sram_data_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_din0[9]  (.DIODE(\SRAMController_ins.sram_data_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0604__X (.DIODE(\SRAMController_ins.sram_data_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[0]  (.DIODE(\SRAMController_ins.sram_data_out[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__A0 (.DIODE(\SRAMController_ins.sram_data_out[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[10]  (.DIODE(\SRAMController_ins.sram_data_out[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__A0 (.DIODE(\SRAMController_ins.sram_data_out[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[12]  (.DIODE(\SRAMController_ins.sram_data_out[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__A0 (.DIODE(\SRAMController_ins.sram_data_out[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[13]  (.DIODE(\SRAMController_ins.sram_data_out[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0965__A0 (.DIODE(\SRAMController_ins.sram_data_out[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[14]  (.DIODE(\SRAMController_ins.sram_data_out[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0967__A0 (.DIODE(\SRAMController_ins.sram_data_out[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[15]  (.DIODE(\SRAMController_ins.sram_data_out[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0969__A0 (.DIODE(\SRAMController_ins.sram_data_out[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[16]  (.DIODE(\SRAMController_ins.sram_data_out[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0971__A0 (.DIODE(\SRAMController_ins.sram_data_out[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[17]  (.DIODE(\SRAMController_ins.sram_data_out[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0973__A0 (.DIODE(\SRAMController_ins.sram_data_out[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[18]  (.DIODE(\SRAMController_ins.sram_data_out[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__A0 (.DIODE(\SRAMController_ins.sram_data_out[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[1]  (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0940__A0 (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[20]  (.DIODE(\SRAMController_ins.sram_data_out[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__A0 (.DIODE(\SRAMController_ins.sram_data_out[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[21]  (.DIODE(\SRAMController_ins.sram_data_out[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__A0 (.DIODE(\SRAMController_ins.sram_data_out[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[22]  (.DIODE(\SRAMController_ins.sram_data_out[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__A0 (.DIODE(\SRAMController_ins.sram_data_out[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[23]  (.DIODE(\SRAMController_ins.sram_data_out[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__A0 (.DIODE(\SRAMController_ins.sram_data_out[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[24]  (.DIODE(\SRAMController_ins.sram_data_out[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0988__A0 (.DIODE(\SRAMController_ins.sram_data_out[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[25]  (.DIODE(\SRAMController_ins.sram_data_out[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__A0 (.DIODE(\SRAMController_ins.sram_data_out[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[26]  (.DIODE(\SRAMController_ins.sram_data_out[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__A0 (.DIODE(\SRAMController_ins.sram_data_out[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[27]  (.DIODE(\SRAMController_ins.sram_data_out[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__A0 (.DIODE(\SRAMController_ins.sram_data_out[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[28]  (.DIODE(\SRAMController_ins.sram_data_out[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__A0 (.DIODE(\SRAMController_ins.sram_data_out[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[29]  (.DIODE(\SRAMController_ins.sram_data_out[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__A0 (.DIODE(\SRAMController_ins.sram_data_out[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[2]  (.DIODE(\SRAMController_ins.sram_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0942__A0 (.DIODE(\SRAMController_ins.sram_data_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[30]  (.DIODE(\SRAMController_ins.sram_data_out[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__A0 (.DIODE(\SRAMController_ins.sram_data_out[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[31]  (.DIODE(\SRAMController_ins.sram_data_out[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1002__A0 (.DIODE(\SRAMController_ins.sram_data_out[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[3]  (.DIODE(\SRAMController_ins.sram_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0944__A0 (.DIODE(\SRAMController_ins.sram_data_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[4]  (.DIODE(\SRAMController_ins.sram_data_out[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0946__A0 (.DIODE(\SRAMController_ins.sram_data_out[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[5]  (.DIODE(\SRAMController_ins.sram_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0948__A0 (.DIODE(\SRAMController_ins.sram_data_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[7]  (.DIODE(\SRAMController_ins.sram_data_out[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0952__A0 (.DIODE(\SRAMController_ins.sram_data_out[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[8]  (.DIODE(\SRAMController_ins.sram_data_out[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0954__A0 (.DIODE(\SRAMController_ins.sram_data_out[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 \ANTENNA_sram_ins_dout0[9]  (.DIODE(\SRAMController_ins.sram_data_out[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0956__A0 (.DIODE(\SRAMController_ins.sram_data_out[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__Q (.DIODE(\SRAMController_ins.sram_tmp[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__A1 (.DIODE(\SRAMController_ins.sram_tmp[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__B2 (.DIODE(\SRAMController_ins.sram_tmp[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1168__Q (.DIODE(\SRAMController_ins.sram_tmp[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__A1 (.DIODE(\SRAMController_ins.sram_tmp[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__B2 (.DIODE(\SRAMController_ins.sram_tmp[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__Q (.DIODE(\SRAMController_ins.sram_tmp[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__A1 (.DIODE(\SRAMController_ins.sram_tmp[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0879__A1 (.DIODE(\SRAMController_ins.sram_tmp[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1170__Q (.DIODE(\SRAMController_ins.sram_tmp[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__A1 (.DIODE(\SRAMController_ins.sram_tmp[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0885__B2 (.DIODE(\SRAMController_ins.sram_tmp[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__Q (.DIODE(\SRAMController_ins.sram_tmp[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0988__A1 (.DIODE(\SRAMController_ins.sram_tmp[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__B2 (.DIODE(\SRAMController_ins.sram_tmp[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1172__Q (.DIODE(\SRAMController_ins.sram_tmp[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__A1 (.DIODE(\SRAMController_ins.sram_tmp[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__A1 (.DIODE(\SRAMController_ins.sram_tmp[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__Q (.DIODE(\SRAMController_ins.sram_tmp[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__A1 (.DIODE(\SRAMController_ins.sram_tmp[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__A1 (.DIODE(\SRAMController_ins.sram_tmp[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1174__Q (.DIODE(\SRAMController_ins.sram_tmp[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__A1 (.DIODE(\SRAMController_ins.sram_tmp[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__A1 (.DIODE(\SRAMController_ins.sram_tmp[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1175__Q (.DIODE(\SRAMController_ins.sram_tmp[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__A1 (.DIODE(\SRAMController_ins.sram_tmp[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0869__A1 (.DIODE(\SRAMController_ins.sram_tmp[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__Q (.DIODE(\SRAMController_ins.sram_tmp[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__A1 (.DIODE(\SRAMController_ins.sram_tmp[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__B2 (.DIODE(\SRAMController_ins.sram_tmp[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__Q (.DIODE(\SRAMController_ins.sram_tmp[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0944__A1 (.DIODE(\SRAMController_ins.sram_tmp[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__A1 (.DIODE(\SRAMController_ins.sram_tmp[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__Q (.DIODE(\SRAMController_ins.sram_tmp[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0946__A1 (.DIODE(\SRAMController_ins.sram_tmp[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__A1 (.DIODE(\SRAMController_ins.sram_tmp[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__Q (.DIODE(\SRAMController_ins.sram_tmp[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0948__A1 (.DIODE(\SRAMController_ins.sram_tmp[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__A1 (.DIODE(\SRAMController_ins.sram_tmp[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__Q (.DIODE(\SRAMController_ins.sram_tmp[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0950__A1 (.DIODE(\SRAMController_ins.sram_tmp[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__A1 (.DIODE(\SRAMController_ins.sram_tmp[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__Q (.DIODE(\SRAMController_ins.sram_tmp[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0952__A1 (.DIODE(\SRAMController_ins.sram_tmp[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0885__A1 (.DIODE(\SRAMController_ins.sram_tmp[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_sram_ins_web0 (.DIODE(\SRAMController_ins.we_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__B (.DIODE(\SRAMController_ins.we_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__B1 (.DIODE(\SRAMController_ins.we_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__B1 (.DIODE(\SRAMController_ins.we_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__B1 (.DIODE(\SRAMController_ins.we_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__B1 (.DIODE(\SRAMController_ins.we_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__A (.DIODE(\SRAMController_ins.we_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0652__X (.DIODE(\SRAMController_ins.we_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0885__A2 (.DIODE(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__A2 (.DIODE(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__A2 (.DIODE(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__A2 (.DIODE(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__A2 (.DIODE(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__A2 (.DIODE(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0855__A2 (.DIODE(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__A2 (.DIODE(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__B1_N (.DIODE(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0557__A1 (.DIODE(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0554__X (.DIODE(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0885__B1 (.DIODE(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0879__A2 (.DIODE(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__B1 (.DIODE(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__B1 (.DIODE(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__B1 (.DIODE(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__B1 (.DIODE(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0855__B1 (.DIODE(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0851__A2 (.DIODE(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__D1 (.DIODE(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0557__A2 (.DIODE(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0555__X (.DIODE(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0884__A2 (.DIODE(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__B1 (.DIODE(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0874__A2 (.DIODE(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0869__A2 (.DIODE(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__A2 (.DIODE(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__A2 (.DIODE(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__A2 (.DIODE(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__B1 (.DIODE(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__B (.DIODE(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0557__A3 (.DIODE(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0556__X (.DIODE(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0648__B (.DIODE(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0646__B (.DIODE(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0644__B (.DIODE(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0642__B (.DIODE(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0640__B (.DIODE(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0638__B (.DIODE(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0636__B (.DIODE(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0615__A (.DIODE(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0594__A (.DIODE(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0583__A (.DIODE(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0582__X (.DIODE(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__A (.DIODE(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__A2 (.DIODE(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__A2 (.DIODE(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__A2 (.DIODE(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__A2 (.DIODE(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0592__B (.DIODE(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0590__B (.DIODE(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0588__B (.DIODE(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0586__B (.DIODE(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0584__B (.DIODE(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0583__X (.DIODE(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0884__B1 (.DIODE(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0879__B1 (.DIODE(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0874__B1 (.DIODE(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0869__B1 (.DIODE(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__B1 (.DIODE(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__B1 (.DIODE(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__B1 (.DIODE(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0851__B1 (.DIODE(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__A2 (.DIODE(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0660__B (.DIODE(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0659__X (.DIODE(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__S (.DIODE(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__S (.DIODE(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__S (.DIODE(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__S (.DIODE(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0667__B1 (.DIODE(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0666__X (.DIODE(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1002__S (.DIODE(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__S (.DIODE(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__A (.DIODE(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0958__A (.DIODE(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0937__A (.DIODE(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__D_N (.DIODE(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__X (.DIODE(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0852__A2 (.DIODE(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0851__X (.DIODE(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0860__A2 (.DIODE(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__X (.DIODE(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0865__B1 (.DIODE(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__X (.DIODE(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__B1 (.DIODE(_0391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__X (.DIODE(_0391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0876__A2 (.DIODE(_0395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__X (.DIODE(_0395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0879__C1 (.DIODE(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__X (.DIODE(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0886__A2 (.DIODE(_0403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0885__X (.DIODE(_0403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0956__S (.DIODE(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0954__S (.DIODE(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0952__S (.DIODE(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0950__S (.DIODE(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0948__S (.DIODE(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0946__S (.DIODE(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0944__S (.DIODE(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0942__S (.DIODE(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0940__S (.DIODE(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__S (.DIODE(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0937__X (.DIODE(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0977__S (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__S (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0973__S (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0971__S (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0969__S (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0967__S (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0965__S (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__S (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0961__S (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__S (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0958__X (.DIODE(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1070__S (.DIODE(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1068__S (.DIODE(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__A (.DIODE(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1026__A (.DIODE(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1005__A (.DIODE(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__X (.DIODE(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout11_X (.DIODE(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0876__A1 (.DIODE(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0856__A1 (.DIODE(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0865__B2 (.DIODE(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__B2 (.DIODE(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0907__B1 (.DIODE(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__A1 (.DIODE(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0660__A_N (.DIODE(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__A_N (.DIODE(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0557__B1 (.DIODE(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0551__B1 (.DIODE(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout16_X (.DIODE(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__RESET_B (.DIODE(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__RESET_B (.DIODE(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__RESET_B (.DIODE(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout14_A (.DIODE(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout15_A (.DIODE(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1214__RESET_B (.DIODE(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1212__RESET_B (.DIODE(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout18_X (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0784__C1 (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout17_A (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__RESET_B (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__RESET_B (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__RESET_B (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1092__RESET_B (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__RESET_B (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout21_X (.DIODE(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__C1 (.DIODE(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__C1 (.DIODE(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0853__C1 (.DIODE(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1182__RESET_B (.DIODE(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__RESET_B (.DIODE(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__RESET_B (.DIODE(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0911__A (.DIODE(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0787__C1 (.DIODE(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0532__A (.DIODE(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0520__B1 (.DIODE(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout23_X (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout21_A (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout22_A (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1166__RESET_B (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1158__RESET_B (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__RESET_B (.DIODE(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout26_X (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0832__A (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0827__C1 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0823__A (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0818__C1 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__C1 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__A (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__0803__C1 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout25_A (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout24_A (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout28_X (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__RESET_B (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout27_A (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__RESET_B (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1172__RESET_B (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1160__RESET_B (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__RESET_B (.DIODE(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout29_X (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout26_A (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout28_A (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout20_A (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout16_A (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout23_A (.DIODE(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload0_A (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__CLK (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__CLK (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__CLK (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1189__CLK (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1192__CLK (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__CLK (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1197__CLK (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1201__CLK (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1202__CLK (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1203__CLK (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1204__CLK (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1205__CLK (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload2_A (.DIODE(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__CLK (.DIODE(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__CLK (.DIODE(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__CLK (.DIODE(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__CLK (.DIODE(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__CLK (.DIODE(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1158__CLK (.DIODE(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1166__CLK (.DIODE(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1199__CLK (.DIODE(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1200__CLK (.DIODE(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_sram_ins_clk0 (.DIODE(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1184__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1190__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1193__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1194__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1196__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1198__CLK (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload7_A (.DIODE(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1109__CLK (.DIODE(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__CLK (.DIODE(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1111__CLK (.DIODE(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__CLK (.DIODE(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload9_A (.DIODE(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__CLK (.DIODE(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__CLK (.DIODE(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1172__CLK (.DIODE(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__CLK (.DIODE(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1174__CLK (.DIODE(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1175__CLK (.DIODE(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload10_A (.DIODE(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1160__CLK (.DIODE(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__CLK (.DIODE(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1168__CLK (.DIODE(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__CLK (.DIODE(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1170__CLK (.DIODE(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1176__CLK (.DIODE(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__CLK (.DIODE(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA__1178__CLK (.DIODE(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\SRAMController_ins.sram_data_out[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\SRAMController_ins.sram_data_out[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\SRAMController_ins.sram_data_out[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\SRAMController_ins.sram_data_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\SRAMController_ins.sram_data_out[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_150 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_378 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_591 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_594 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_597 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_603 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_638 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_651 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_657 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_660 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_667 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_677 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_688 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_769 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_772 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_797 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_803 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_843 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_855 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_981 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1013 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1025 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1059 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1016 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1038 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1050 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1062 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1074 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1086 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_115 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1038 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1018 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1022 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1055 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1067 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1079 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1027 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1016 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1047 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1059 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1071 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1083 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1018 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1025 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1051 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_108 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1036 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_132 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1046 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1058 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1066 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_106 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1016 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1030 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1038 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1016 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1046 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1058 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1066 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1016 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1025 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1037 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_136 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1024 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1036 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1048 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1060 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1018 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1030 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1066 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_118 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1027 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1039 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_144 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1033 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1045 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1057 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_128 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1038 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1016 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1044 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1056 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1019 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1031 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1039 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1019 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1031 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1043 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1055 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1067 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_127 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1019 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1031 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1039 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1043 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1055 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1067 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1018 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1030 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1038 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1019 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1031 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1039 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_172 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1025 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1031 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1039 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1031 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1043 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1055 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1067 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1027 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1039 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_170 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_155 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_166 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1019 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1031 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1039 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1019 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1031 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1043 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1055 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1067 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1042 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1054 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1066 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1078 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1016 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1028 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1040 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1052 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1070 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_256 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_268 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_281 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_293 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_337 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_395 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_407 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_449 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_494 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_501 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_505 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_517 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_561 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_573 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_600 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_619 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_631 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_645 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_657 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_673 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_685 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_701 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_713 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_729 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_741 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_753 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_765 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_782 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_785 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_797 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_809 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_813 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_825 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_837 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_841 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_853 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_865 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_869 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_881 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_893 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_897 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_909 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_921 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_925 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_937 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_953 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_965 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_977 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_981 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_993 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_369 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_462 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_471 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_539 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_568 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_621 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_634 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_648 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_660 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_673 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_685 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_697 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_709 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_713 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_717 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_738 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_746 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_751 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_763 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_780 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_785 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_797 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_809 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_821 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_833 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_841 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_853 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_865 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_877 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_889 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_897 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_909 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_921 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_933 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_945 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_953 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_965 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_977 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_989 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1033 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1045 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_448 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_459 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_511 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_519 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_535 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_578 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_593 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_596 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_607 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_626 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_648 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_775 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_787 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_799 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_813 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_825 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_837 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_849 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_861 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_869 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_881 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_893 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_905 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_917 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_925 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_937 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_949 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_961 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_973 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_981 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_993 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1005 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1017 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1029 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1061 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1073 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_430 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_507 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_513 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_541 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_547 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_583 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_591 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_646 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_652 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_768 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_780 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_785 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_797 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_809 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_821 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_833 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_841 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_853 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_865 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_877 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_889 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_897 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_909 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_921 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_933 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_945 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_953 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_965 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_977 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_989 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1033 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1045 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_225 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_509 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_541 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_546 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_572 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_576 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_591 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_599 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_657 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_678 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_709 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_719 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_731 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_775 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_787 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_799 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_813 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_825 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_837 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_849 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_861 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_869 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_881 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_893 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_905 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_917 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_925 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_937 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_949 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_961 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_973 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_981 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_993 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1005 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1017 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1029 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1061 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1073 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_197 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_253 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_289 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_367 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_467 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_471 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_483 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_495 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_535 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_603 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_649 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_666 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_681 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_705 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_717 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_745 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_762 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_774 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_782 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_785 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_797 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_809 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_821 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_833 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_841 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_853 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_865 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_877 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_889 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_897 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_909 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_921 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_933 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_945 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_953 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_965 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_977 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_989 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1033 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1045 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_157 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_200 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_220 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_374 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_404 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_460 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_472 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_545 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_564 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_572 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_582 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_607 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_619 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_648 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_654 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_677 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_701 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_713 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_725 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_737 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_757 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_769 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_781 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_793 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_805 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_813 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_825 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_837 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_849 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_861 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_869 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_881 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_893 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_905 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_917 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_925 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_937 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_949 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_961 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_973 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_981 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_993 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1005 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1017 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1029 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1061 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1073 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_187 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_400 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_412 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_424 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_436 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_577 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_597 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_604 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_611 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_651 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_681 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_704 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_760 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_772 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_785 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_797 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_809 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_821 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_833 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_841 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_853 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_865 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_877 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_889 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_897 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_909 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_921 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_933 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_945 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_953 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_965 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_977 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_989 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1033 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1045 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_227 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_239 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_565 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_575 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_742 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_754 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_757 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_769 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_781 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_793 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_805 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_813 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_825 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_837 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_849 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_861 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_869 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_881 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_893 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_905 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_917 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_925 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_937 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_949 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_961 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_973 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_981 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_993 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1005 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1017 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1029 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1061 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1073 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_411 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_423 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_435 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_579 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_705 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_737 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_770 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_782 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_785 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_797 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_809 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_821 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_833 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_841 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_853 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_865 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_877 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_889 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_897 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_909 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_921 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_933 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_945 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_953 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_965 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_977 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_989 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1033 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1045 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_154 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_225 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_237 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_283 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_324 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_337 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_349 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_449 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_461 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_501 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_505 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_517 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_561 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_573 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_632 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_658 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_704 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_716 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_729 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_744 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_769 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_781 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_785 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_797 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_809 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_813 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_825 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_837 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_841 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_853 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_865 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_869 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_881 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_893 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_897 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_909 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_921 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_925 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_937 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_953 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_965 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_977 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_981 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_993 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1009 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1021 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1037 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1049 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1065 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1077 (.VPWR(VDPWR),
    .VGND(VGND),
    .VPB(VDPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VDPWR),
    .VPWR(VDPWR));
 assign uio_oe[0] = net35;
 assign uio_oe[1] = net36;
 assign uio_oe[2] = net37;
 assign uio_oe[3] = net38;
 assign uio_oe[4] = net56;
 assign uio_oe[5] = net39;
 assign uio_oe[6] = net40;
 assign uio_oe[7] = net41;
 assign uio_out[0] = net42;
 assign uio_out[1] = net43;
 assign uio_out[2] = net44;
 assign uio_out[3] = net45;
 assign uio_out[5] = net46;
 assign uio_out[6] = net47;
 assign uio_out[7] = net48;
 assign uo_out[0] = net49;
 assign uo_out[1] = net50;
 assign uo_out[2] = net51;
 assign uo_out[3] = net52;
 assign uo_out[4] = net53;
 assign uo_out[5] = net54;
endmodule
